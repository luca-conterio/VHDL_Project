----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 12.12.2017 17:48:44
-- Design Name: 
-- Module Name: FSM_testbench - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
 
entity project_tb is
end project_tb;


architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 15 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst		    : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		    : std_logic := '0';
signal   mem_o_data,mem_i_data		: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		: std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (2 => "10110000", 3 => "10100110", 4 => "10111001", 6 => "00001011", 7 => "10001101", 8 => "10111101", 9 => "01101110", 10 => "10110010", 11 => "01101011", 12 => "11110101", 14 => "10011110", 15 => "00101111", 16 => "01011001", 17 => "01100001", 18 => "00100011", 21 => "01110000", 22 => "00010110", 23 => "01011100", 24 => "01100011", 25 => "10101111", 26 => "11010000", 27 => "10000110", 28 => "10001100", 29 => "11111111", 30 => "00111100", 31 => "11001111", 32 => "10010000", 35 => "01011100", 36 => "00001010", 37 => "00100000", 38 => "10000100", 39 => "01010111", 40 => "10100001", 41 => "00111101", 42 => "10110010", 43 => "10010101", 44 => "10111100", 45 => "01001000", 46 => "00011010", 48 => "11010100", 53 => "11101110", 54 => "00110011", 56 => "11001011", 57 => "00110000", 60 => "11110111", 63 => "00011011", 65 => "10000010", 66 => "11001100", 67 => "01110111", 69 => "00111101", 70 => "10011111", 71 => "10110001", 73 => "10110011", 76 => "10101101", 77 => "11000001", 78 => "11111100", 79 => "00100101", 82 => "10001011", 85 => "01001111", 87 => "11001011", 88 => "10111010", 89 => "00000111", 90 => "11101101", 91 => "10110010", 92 => "01111000", 94 => "00010010", 95 => "01111001", 99 => "10011010", 100 => "10100001", 101 => "00011110", 102 => "00111100", 107 => "11010101", 110 => "10110001", 111 => "01100100", 112 => "00101010", 113 => "11001001", 114 => "11001101", 117 => "01001011", 120 => "01101011", 121 => "10010010", 122 => "00110110", 123 => "00111010", 125 => "10110000", 126 => "11001101", 128 => "10111100", 129 => "01011101", 130 => "10111101", 131 => "01010111", 132 => "01111010", 133 => "01010001", 135 => "00110101", 136 => "01000111", 138 => "11001000", 139 => "11010001", 140 => "11111110", 144 => "01111010", 145 => "10010011", 146 => "11001001", 147 => "00101001", 148 => "00001011", 149 => "00101001", 150 => "01110011", 151 => "10100000", 153 => "10111000", 154 => "11001000", 155 => "10110100", 157 => "11000001", 158 => "11110110", 160 => "00101011", 161 => "01101100", 163 => "00011101", 164 => "00000011", 165 => "10110100", 166 => "10010101", 167 => "01110111", 168 => "11110001", 169 => "01011110", 171 => "00100111", 172 => "10000001", 175 => "00001011", 177 => "10111100", 179 => "10000000", 180 => "10000101", 181 => "10110110", 182 => "00100100", 184 => "11010101", 186 => "01000011", 189 => "01110001", 190 => "10111100", 191 => "11111100", 192 => "00100111", 193 => "00011111", 195 => "01010100", 197 => "10111110", 198 => "11011100", 199 => "10110101", 200 => "10011011", 201 => "11011100", 203 => "00000011", 205 => "00101111", 206 => "10011100", 208 => "10100010", 210 => "10011110", 211 => "00011010", 212 => "00000101", 215 => "10110101", 216 => "10001100", 217 => "00001100", 218 => "00011000", 219 => "10101010", 220 => "11111111", 221 => "00011100", 223 => "10001100", 224 => "00010101", 225 => "01101101", 226 => "11110110", 228 => "00101110", 229 => "11100110", 230 => "10110011", 232 => "10000000", 234 => "10010001", 236 => "11101101", 237 => "11100001", 240 => "00011011", 242 => "10111110", 243 => "10010111", 244 => "11001111", 245 => "11010100", 246 => "01010000", 248 => "00101011", 249 => "10000100", 250 => "00011111", 251 => "11001111", 252 => "10011100", 254 => "11111011", 255 => "10110111", 256 => "11110011", 258 => "01100011", 259 => "11100110", 260 => "00001000", 261 => "10000100", 262 => "00110010", 263 => "00011110", 264 => "01010101", 265 => "11011001", 266 => "10010110", 267 => "11111001", 268 => "11011110", 270 => "10101001", 271 => "00001110", 273 => "10100011", 274 => "10101110", 275 => "01000011", 276 => "10000101", 280 => "11111100", 282 => "01110111", 284 => "11110110", 285 => "00010011", 288 => "10110000", 289 => "11000110", 290 => "10101111", 292 => "00111010", 293 => "01100111", 294 => "11011000", 296 => "01011111", 298 => "11001111", 300 => "11011101", 301 => "10111100", 302 => "10111000", 303 => "10001101", 305 => "10000100", 306 => "11001100", 307 => "11010001", 309 => "00001101", 310 => "10001011", 311 => "01011110", 312 => "11101111", 313 => "01000100", 316 => "01010111", 317 => "11101111", 318 => "00100111", 319 => "01001011", 320 => "10101101", 321 => "01000000", 322 => "11011110", 323 => "00111101", 325 => "01010001", 326 => "10000110", 327 => "01001001", 328 => "10111011", 330 => "11001101", 331 => "10100101", 332 => "00101100", 333 => "00100011", 334 => "11001101", 336 => "01000011", 337 => "10110101", 338 => "00011100", 339 => "01010100", 340 => "00100111", 341 => "00110111", 342 => "10101000", 343 => "00101010", 344 => "11110111", 346 => "00011000", 347 => "00111110", 348 => "10001011", 351 => "01010110", 352 => "00110101", 353 => "00100101", 354 => "11010111", 355 => "10100110", 356 => "01010000", 357 => "10111110", 358 => "10000111", 359 => "00000011", 360 => "00111000", 361 => "10111110", 362 => "11010110", 363 => "00110100", 364 => "01100111", 365 => "11110101", 367 => "10000001", 368 => "01100111", 371 => "01101110", 373 => "01100001", 374 => "01010011", 375 => "11110011", 377 => "00111101", 378 => "11010111", 379 => "01011000", 380 => "10111001", 381 => "00011111", 383 => "00110001", 384 => "11111010", 386 => "10001111", 387 => "11110000", 388 => "00101001", 389 => "01111001", 390 => "11001010", 391 => "10110001", 392 => "00011010", 397 => "10110000", 399 => "00100010", 400 => "00111010", 401 => "00011101", 402 => "10011010", 403 => "00111110", 404 => "00011000", 405 => "11111010", 406 => "00001100", 407 => "00000001", 408 => "00111010", 409 => "10001010", 412 => "01011000", 413 => "00100001", 415 => "11001111", 416 => "11010101", 419 => "11000011", 420 => "11010110", 421 => "11111111", 422 => "01110011", 423 => "11110011", 424 => "10000100", 425 => "01000010", 426 => "01010000", 427 => "01001011", 428 => "11110101", 429 => "01111011", 430 => "01110011", 431 => "10110000", 432 => "00110011", 433 => "11101111", 434 => "01111101", 435 => "11010101", 436 => "11010100", 437 => "11100100", 438 => "00011110", 441 => "10010000", 442 => "00011001", 443 => "11011000", 444 => "01001110", 445 => "11101011", 446 => "00100101", 447 => "11110010", 451 => "01110000", 452 => "10000101", 454 => "11001101", 457 => "10101000", 459 => "10000001", 461 => "00010000", 462 => "00111111", 463 => "10000100", 464 => "00100100", 465 => "01111110", 466 => "10100101", 467 => "00111110", 468 => "11110101", 471 => "11000111", 472 => "01110001", 473 => "10100111", 474 => "01100110", 475 => "01000110", 477 => "00011011", 478 => "10001001", 479 => "01100011", 480 => "10000001", 482 => "00001111", 484 => "11001000", 485 => "11100010", 487 => "00001100", 488 => "01101111", 489 => "11011000", 490 => "00011011", 491 => "01110001", 492 => "11010111", 493 => "11001010", 494 => "11000010", 496 => "11001001", 498 => "10011001", 499 => "11100101", 500 => "11110100", 501 => "11010010", 502 => "01111011", 503 => "00001001", 504 => "11000011", 505 => "00011101", 509 => "10010010", 510 => "00101100", 512 => "11111001", 513 => "10110001", 514 => "10110111", 515 => "11110101", 516 => "01100101", 518 => "11100010", 519 => "10101111", 520 => "10011101", 521 => "00101000", 522 => "11001011", 523 => "10110001", 524 => "10111111", 525 => "11000011", 527 => "10010001", 528 => "11010010", 529 => "00100010", 530 => "01101011", 531 => "10001001", 532 => "11011011", 533 => "01001000", 534 => "10101101", 535 => "10100101", 536 => "10000100", 537 => "00011001", 538 => "11010000", 540 => "01111100", 541 => "00110000", 542 => "11001101", 543 => "10111111", 545 => "11100110", 546 => "10110101", 548 => "11011001", 551 => "11011101", 552 => "00110001", 554 => "01011111", 555 => "00000100", 556 => "10011010", 557 => "10110110", 558 => "11100111", 560 => "10000110", 561 => "10101100", 563 => "10011110", 564 => "10010001", 565 => "10000011", 566 => "11110111", 567 => "00000010", 568 => "11001100", 569 => "11010000", 570 => "10110001", 571 => "00100111", 572 => "10110010", 573 => "11110000", 575 => "10110010", 576 => "01100010", 578 => "11100100", 579 => "10100011", 580 => "10110110", 583 => "00100011", 584 => "01011000", 585 => "10100000", 587 => "01101101", 588 => "01001011", 590 => "00000011", 591 => "10001011", 592 => "00001101", 594 => "00010100", 595 => "01110011", 597 => "01010001", 598 => "11111101", 599 => "11011100", 600 => "00001111", 601 => "00101001", 603 => "11101110", 604 => "00000011", 605 => "10011110", 606 => "01100101", 608 => "00001111", 609 => "01101101", 610 => "11110010", 612 => "00111011", 613 => "11110001", 614 => "00111101", 615 => "11000110", 616 => "00101000", 617 => "11011001", 622 => "10111001", 623 => "00111000", 624 => "01011001", 630 => "11011101", 632 => "11000011", 633 => "00010001", 637 => "00001011", 638 => "10000001", 639 => "10100100", 640 => "10111011", 641 => "00110000", 642 => "11011000", 643 => "10110000", 644 => "10000110", 645 => "01001101", 646 => "11111100", 647 => "01001101", 649 => "11110000", 650 => "01011110", 651 => "00010011", 652 => "10101011", 653 => "11100110", 654 => "11100001", 655 => "01000011", 657 => "01001000", 660 => "10010010", 663 => "00111110", 664 => "10000001", 666 => "00101100", 667 => "01001011", 669 => "00110010", 670 => "00101001", 671 => "11001101", 672 => "11000000", 673 => "01001100", 674 => "00001000", 675 => "11000110", 676 => "11001010", 677 => "11001101", 678 => "10100100", 682 => "00001111", 683 => "01011111", 685 => "11000011", 686 => "11011001", 687 => "10010111", 688 => "11000000", 691 => "10011100", 692 => "11011001", 693 => "11100010", 694 => "00111111", 696 => "11100001", 697 => "00100001", 699 => "10111010", 700 => "11010001", 701 => "10000010", 702 => "01010110", 704 => "00000110", 707 => "01100101", 710 => "01101111", 711 => "11011101", 712 => "11110010", 713 => "00111010", 714 => "10011110", 715 => "00110001", 717 => "11011110", 720 => "00011010", 724 => "00111111", 725 => "01101010", 726 => "11001100", 727 => "00010011", 728 => "10010101", 730 => "10010110", 731 => "11011001", 732 => "11001111", 733 => "00101110", 735 => "10101100", 736 => "10010101", 737 => "11001010", 738 => "01001001", 739 => "00011110", 740 => "10110011", 741 => "00010000", 742 => "01101010", 743 => "10110011", 744 => "00110101", 747 => "11111011", 748 => "11100101", 751 => "00101010", 752 => "10011001", 753 => "00110110", 754 => "10010001", 755 => "01000110", 757 => "11011110", 758 => "11101100", 759 => "01011110", 760 => "01101100", 761 => "01001111", 762 => "00110001", 763 => "10111101", 764 => "11001010", 765 => "10001000", 766 => "11011011", 769 => "01000100", 770 => "00111110", 771 => "10001100", 772 => "01100011", 774 => "10001000", 775 => "10010100", 777 => "11101110", 778 => "10011001", 779 => "00111110", 780 => "11110100", 784 => "01000001", 785 => "10110111", 786 => "11010101", 788 => "01011011", 789 => "01000110", 791 => "00010101", 793 => "10001101", 794 => "01110101", 795 => "11101111", 796 => "11010001", 798 => "00001011", 799 => "01111110", 800 => "11110100", 801 => "11100110", 802 => "00100001", 803 => "01101010", 804 => "10010010", 806 => "11111111", 807 => "11000100", 808 => "11101000", 809 => "00011100", 810 => "10101001", 812 => "00110011", 813 => "10010000", 814 => "01000101", 815 => "10010101", 816 => "11011001", 817 => "00001110", 818 => "01101110", 819 => "11111011", 820 => "01110100", 821 => "10000100", 822 => "10011101", 823 => "01010011", 824 => "10001101", 825 => "10011101", 826 => "00001001", 827 => "10000010", 829 => "11011011", 830 => "00011011", 831 => "01001101", 832 => "00010011", 833 => "11110111", 836 => "11100101", 837 => "01101010", 838 => "00110111", 839 => "00111011", 844 => "00111010", 845 => "10101000", 848 => "10101001", 849 => "01010100", 855 => "11011101", 856 => "01000000", 857 => "11001010", 858 => "01111010", 860 => "01111000", 861 => "00000110", 862 => "00110011", 864 => "11011011", 865 => "00010001", 866 => "11100110", 867 => "10101111", 869 => "10001111", 870 => "01010011", 872 => "01101111", 873 => "00111001", 874 => "11110100", 876 => "00100110", 877 => "10010100", 879 => "00001011", 880 => "11101100", 882 => "10101101", 883 => "00110011", 884 => "00101111", 885 => "01100011", 886 => "11000010", 887 => "10100001", 888 => "00110111", 889 => "11001001", 890 => "01010110", 892 => "01010001", 894 => "10110011", 895 => "11101001", 896 => "00011010", 898 => "01110000", 900 => "01110110", 901 => "01110001", 902 => "10110001", 904 => "00010111", 905 => "10000101", 906 => "10011100", 908 => "00100111", 909 => "01001101", 910 => "01011011", 911 => "00010001", 912 => "01110111", 913 => "01011111", 915 => "10101011", 916 => "01110001", 917 => "11001000", 918 => "11001001", 919 => "00111010", 921 => "00100010", 924 => "00100011", 925 => "11101010", 927 => "00011111", 929 => "01000111", 930 => "11000000", 932 => "00111001", 933 => "10111110", 934 => "11001101", 935 => "10110100", 936 => "10000100", 937 => "11011001", 938 => "10011011", 939 => "00011100", 941 => "10000101", 942 => "01011111", 945 => "10010010", 946 => "01001000", 947 => "10001100", 948 => "11101000", 949 => "01010110", 950 => "01100100", 951 => "11111100", 952 => "10011000", 953 => "10101001", 955 => "00100001", 956 => "01100110", 957 => "01001011", 958 => "11101010", 960 => "10101000", 961 => "01101100", 962 => "10110100", 963 => "01001001", 964 => "01011111", 965 => "00010010", 966 => "01010000", 967 => "01011010", 969 => "00111011", 970 => "10010001", 971 => "11010010", 972 => "01010001", 973 => "00111001", 975 => "11010010", 976 => "11110100", 977 => "11011001", 978 => "11110010", 980 => "10010011", 982 => "10111101", 983 => "01011110", 984 => "00000110", 986 => "01010101", 987 => "11010100", 988 => "11100011", 989 => "11000100", 990 => "01100111", 992 => "10010100", 993 => "11011011", 994 => "11111010", 995 => "00110001", 996 => "11000001", 997 => "11101001", 998 => "11111100", 999 => "00110100", 1000 => "01000010", 1001 => "01110011", 1002 => "11000101", 1003 => "01001000", 1004 => "11101110", 1005 => "11001111", 1006 => "10101000", 1007 => "00011111", 1008 => "10001101", 1009 => "00001011", 1011 => "11011010", 1012 => "11101111", 1013 => "11110110", 1014 => "01000001", 1015 => "11010100", 1016 => "11010110", 1017 => "11000011", 1018 => "11100111", 1020 => "10011111", 1021 => "10000101", 1023 => "01011110", 1024 => "11011100", 1025 => "10100000", 1026 => "10000011", 1027 => "10011010", 1030 => "00100110", 1031 => "01010111", 1032 => "11000110", 1033 => "11010101", 1035 => "11101000", 1036 => "00001000", 1037 => "10111111", 1038 => "00010100", 1039 => "00011111", 1040 => "01010111", 1042 => "10011010", 1044 => "11001110", 1045 => "10001100", 1047 => "10000001", 1051 => "10011110", 1052 => "10111000", 1055 => "10000101", 1056 => "11011010", 1057 => "10101000", 1058 => "11000000", 1059 => "00100111", 1060 => "11000011", 1061 => "01111011", 1063 => "01101001", 1064 => "01011110", 1065 => "10001011", 1067 => "10110100", 1068 => "10101101", 1069 => "11000000", 1070 => "11010001", 1071 => "00101010", 1072 => "01010111", 1075 => "10110111", 1077 => "10110111", 1078 => "10110010", 1079 => "11001110", 1080 => "11010000", 1083 => "01011001", 1086 => "00010111", 1087 => "01010001", 1088 => "10110101", 1090 => "00100111", 1091 => "00010110", 1093 => "10111110", 1094 => "11011101", 1095 => "10011001", 1097 => "00000011", 1100 => "00111010", 1101 => "10110011", 1103 => "00010101", 1104 => "00001001", 1105 => "00010110", 1106 => "11100001", 1107 => "10111010", 1108 => "11110100", 1110 => "10111101", 1112 => "10010010", 1113 => "00011011", 1114 => "10110101", 1115 => "11101100", 1116 => "11000111", 1117 => "10011000", 1119 => "10001110", 1120 => "00111111", 1121 => "00110111", 1122 => "10010100", 1123 => "10100010", 1124 => "10011110", 1127 => "01010011", 1128 => "01011001", 1129 => "00011101", 1130 => "00001001", 1131 => "00101100", 1133 => "01001010", 1134 => "01101011", 1135 => "10010100", 1136 => "10110001", 1138 => "11111001", 1140 => "10100001", 1141 => "11111011", 1142 => "00000111", 1144 => "10101010", 1145 => "10010101", 1147 => "01001100", 1152 => "01110100", 1153 => "01001101", 1155 => "00100101", 1156 => "00000011", 1157 => "01110100", 1158 => "10001101", 1161 => "10010001", 1162 => "11100111", 1163 => "11000011", 1164 => "10011110", 1165 => "11001110", 1166 => "01101010", 1167 => "01001000", 1168 => "00111101", 1169 => "01010011", 1170 => "11011011", 1171 => "00010011", 1172 => "01101010", 1174 => "01010111", 1176 => "01111010", 1177 => "00101010", 1178 => "00001011", 1179 => "01101111", 1180 => "00000011", 1181 => "00111111", 1182 => "01100100", 1183 => "10101101", 1184 => "10010010", 1185 => "01101001", 1186 => "11101001", 1187 => "01111001", 1188 => "10011001", 1190 => "10011011", 1191 => "10010101", 1192 => "01011011", 1193 => "11100011", 1195 => "10010011", 1197 => "11101001", 1198 => "11011110", 1199 => "01011101", 1200 => "10000010", 1201 => "11100100", 1202 => "01001010", 1203 => "01111101", 1205 => "00100100", 1206 => "01110100", 1207 => "11111000", 1208 => "10101001", 1209 => "01111110", 1210 => "11001100", 1212 => "00001010", 1213 => "00001100", 1214 => "10101000", 1217 => "01000010", 1219 => "01110111", 1220 => "11011010", 1221 => "00111000", 1222 => "01011001", 1223 => "00110001", 1224 => "01000100", 1225 => "01011001", 1226 => "10111101", 1227 => "10000010", 1228 => "01011110", 1229 => "10110010", 1231 => "10110011", 1232 => "00001110", 1233 => "00100101", 1234 => "01100101", 1235 => "00011101", 1236 => "01011111", 1237 => "01110111", 1238 => "10010010", 1239 => "00101111", 1240 => "00011101", 1242 => "11100001", 1243 => "10110000", 1244 => "01100011", 1245 => "11011111", 1247 => "01101001", 1248 => "10011110", 1250 => "00001000", 1251 => "10111101", 1253 => "10100000", 1255 => "00011011", 1256 => "00010111", 1257 => "11010100", 1260 => "10100111", 1262 => "11000100", 1263 => "10010101", 1264 => "01110011", 1265 => "01100000", 1266 => "00010101", 1267 => "01111110", 1268 => "01000011", 1269 => "11101101", 1270 => "11011100", 1271 => "00111101", 1272 => "11010110", 1273 => "11111111", 1274 => "10000110", 1275 => "01001000", 1276 => "10010110", 1277 => "01101110", 1278 => "00001101", 1279 => "01111110", 1280 => "01101000", 1281 => "01101111", 1282 => "01011111", 1284 => "11100001", 1285 => "10101100", 1287 => "01010100", 1288 => "00011010", 1289 => "01000010", 1290 => "00010010", 1291 => "11011100", 1292 => "10100001", 1293 => "10000001", 1294 => "11000010", 1295 => "10100111", 1297 => "11101011", 1298 => "00101111", 1300 => "01111000", 1301 => "11000010", 1302 => "11010000", 1303 => "01000010", 1306 => "01100010", 1308 => "00011111", 1309 => "11001101", 1310 => "00001100", 1311 => "11010011", 1312 => "10110111", 1313 => "00110100", 1314 => "00101101", 1315 => "11011101", 1316 => "01000001", 1317 => "10110111", 1318 => "00000100", 1319 => "10110101", 1320 => "11111010", 1321 => "10010110", 1322 => "11101000", 1323 => "10010100", 1324 => "01011100", 1325 => "11101111", 1327 => "11110010", 1328 => "10110000", 1330 => "00011000", 1333 => "11110011", 1334 => "00001111", 1335 => "11111110", 1337 => "11101001", 1338 => "11010001", 1339 => "00111101", 1342 => "10000001", 1343 => "00101100", 1344 => "10011101", 1345 => "00001000", 1346 => "10010110", 1348 => "11101001", 1350 => "01101010", 1351 => "00001111", 1352 => "11110001", 1353 => "00010011", 1354 => "00101011", 1355 => "11111000", 1356 => "10010000", 1357 => "11001000", 1358 => "10011100", 1359 => "01010110", 1360 => "10100101", 1361 => "01011011", 1362 => "10011001", 1365 => "11100110", 1366 => "00100011", 1367 => "00110011", 1368 => "10001001", 1369 => "10011111", 1370 => "11111111", 1373 => "01100111", 1374 => "01100001", 1375 => "11110011", 1378 => "00011000", 1381 => "01111011", 1383 => "00011001", 1384 => "10001100", 1385 => "01101010", 1387 => "10100000", 1388 => "01100111", 1389 => "00110001", 1390 => "11101000", 1392 => "11011001", 1393 => "01010010", 1394 => "00011000", 1395 => "00010110", 1396 => "11100111", 1397 => "11000000", 1398 => "11110011", 1399 => "11110111", 1400 => "10010011", 1402 => "10110001", 1404 => "01000111", 1406 => "01010100", 1408 => "01100011", 1409 => "10100111", 1410 => "11111001", 1411 => "10001110", 1412 => "10101001", 1414 => "00001011", 1415 => "01101110", 1417 => "11111011", 1418 => "11101011", 1419 => "11000001", 1420 => "11111011", 1421 => "00101011", 1422 => "10110001", 1423 => "01100111", 1424 => "01011111", 1425 => "11100101", 1426 => "11101100", 1428 => "10100100", 1430 => "00111111", 1431 => "11000111", 1432 => "01011110", 1433 => "01010100", 1434 => "01101100", 1436 => "00111101", 1437 => "01100011", 1439 => "00111011", 1440 => "11001110", 1441 => "10110011", 1443 => "10011001", 1446 => "01001001", 1447 => "11001000", 1449 => "10000001", 1451 => "11000000", 1452 => "01111010", 1453 => "01111101", 1454 => "01000111", 1456 => "10111001", 1458 => "10111110", 1459 => "11111011", 1460 => "01000001", 1463 => "01101000", 1464 => "10110010", 1465 => "11101011", 1466 => "00110010", 1467 => "00100000", 1468 => "01100011", 1471 => "01101000", 1472 => "10011011", 1473 => "01110011", 1474 => "10111000", 1475 => "01111011", 1477 => "11011110", 1478 => "01101001", 1479 => "11001100", 1480 => "01100111", 1483 => "10001010", 1484 => "10001001", 1485 => "11010000", 1486 => "10110011", 1487 => "01111001", 1488 => "10000111", 1489 => "11100010", 1491 => "11111101", 1492 => "10111000", 1493 => "01110011", 1495 => "01011101", 1496 => "01111011", 1498 => "11010111", 1499 => "01010100", 1500 => "11101000", 1501 => "10010110", 1502 => "00001111", 1503 => "10110110", 1504 => "01001010", 1505 => "01111001", 1506 => "10011010", 1507 => "00100101", 1508 => "00100101", 1509 => "11001101", 1510 => "00001010", 1511 => "00000010", 1512 => "11011001", 1513 => "10010010", 1514 => "00001101", 1515 => "11000100", 1516 => "10001011", 1517 => "01011000", 1518 => "10101001", 1519 => "11110011", 1522 => "00101111", 1523 => "00100010", 1524 => "01001010", 1526 => "00101001", 1527 => "00001001", 1528 => "10110111", 1531 => "01111111", 1533 => "10010000", 1536 => "01000011", 1537 => "11111100", 1539 => "01000011", 1540 => "01101000", 1542 => "00101100", 1543 => "11010010", 1544 => "01001111", 1545 => "00010001", 1546 => "01101011", 1547 => "11111111", 1548 => "01001101", 1549 => "10000001", 1550 => "00101100", 1552 => "10110011", 1553 => "01011101", 1555 => "00111111", 1556 => "11100011", 1557 => "11010100", 1559 => "10111110", 1560 => "10100001", 1561 => "11101001", 1566 => "11010001", 1567 => "11000101", 1568 => "01010100", 1569 => "01001010", 1570 => "11000101", 1571 => "00100001", 1572 => "00001010", 1573 => "01100011", 1574 => "10111000", 1579 => "10101110", 1580 => "01011110", 1581 => "10111001", 1582 => "10011000", 1584 => "11000011", 1585 => "10101011", 1586 => "01001011", 1590 => "10001001", 1591 => "01000110", 1592 => "00000111", 1593 => "01100001", 1594 => "10101100", 1596 => "10110101", 1597 => "00010101", 1601 => "01101100", 1602 => "11101101", 1603 => "11100010", 1604 => "10111100", 1605 => "10100000", 1606 => "10011101", 1608 => "01111001", 1609 => "11110110", 1610 => "10010111", 1611 => "10000100", 1612 => "10011010", 1613 => "10100001", 1615 => "11111101", 1616 => "11110001", 1617 => "01110101", 1618 => "10011011", 1620 => "00101111", 1621 => "00111111", 1622 => "10110000", 1623 => "11000010", 1625 => "10111110", 1626 => "11000100", 1627 => "01110000", 1628 => "00101111", 1629 => "11111001", 1630 => "00111101", 1632 => "11010001", 1634 => "11100011", 1635 => "10111101", 1637 => "11110000", 1638 => "10110000", 1640 => "00111010", 1641 => "01111110", 1642 => "01111110", 1643 => "10000001", 1644 => "11111011", 1645 => "11000000", 1646 => "10011011", 1647 => "10000011", 1648 => "10110011", 1649 => "00111110", 1651 => "01100100", 1652 => "00111111", 1654 => "01101111", 1656 => "10110000", 1657 => "11111000", 1658 => "01101101", 1659 => "11100000", 1660 => "10010100", 1661 => "00001001", 1662 => "10101010", 1663 => "01101111", 1664 => "11011100", 1665 => "10000111", 1666 => "01011011", 1667 => "10100001", 1668 => "00000101", 1669 => "10011000", 1671 => "00000100", 1672 => "00011000", 1673 => "10011011", 1674 => "01101011", 1675 => "01111001", 1676 => "10111010", 1677 => "11010011", 1678 => "00111011", 1679 => "00000011", 1680 => "10111100", 1681 => "01010101", 1682 => "10110001", 1683 => "00101001", 1684 => "00111001", 1685 => "10110000", 1686 => "01001111", 1687 => "01001001", 1690 => "11111100", 1694 => "10011101", 1695 => "01010011", 1697 => "11000100", 1698 => "10100000", 1699 => "01010101", 1700 => "01100100", 1701 => "00101111", 1703 => "00010110", 1705 => "10110010", 1706 => "01100100", 1707 => "00111000", 1708 => "01110111", 1709 => "11001001", 1711 => "01011000", 1712 => "00001111", 1713 => "10001000", 1715 => "00000010", 1716 => "00011011", 1717 => "01110111", 1718 => "11111000", 1719 => "00111010", 1720 => "11100001", 1722 => "11110110", 1723 => "00100111", 1725 => "10111000", 1728 => "11001100", 1731 => "11101111", 1732 => "00101001", 1736 => "01110101", 1737 => "01001000", 1738 => "00000100", 1739 => "00011011", 1741 => "11110001", 1742 => "01101010", 1744 => "00000011", 1745 => "00101101", 1746 => "11101011", 1750 => "00010110", 1751 => "10010000", 1752 => "10011101", 1754 => "00011011", 1759 => "01011000", 1760 => "11001100", 1761 => "00110011", 1762 => "01001001", 1764 => "11000110", 1765 => "10101101", 1767 => "01000110", 1768 => "01110010", 1769 => "00100001", 1770 => "01000000", 1771 => "11010000", 1772 => "10100100", 1773 => "11011001", 1774 => "01110111", 1777 => "01101110", 1778 => "01011101", 1781 => "11011001", 1782 => "10110101", 1783 => "10101010", 1785 => "00001111", 1786 => "00111010", 1787 => "00101100", 1789 => "10000111", 1790 => "01001000", 1791 => "01010010", 1792 => "11000111", 1793 => "10001100", 1794 => "11100111", 1795 => "00100110", 1796 => "10101000", 1799 => "01110010", 1800 => "11011000", 1801 => "00100000", 1802 => "10010000", 1803 => "00010110", 1804 => "10011001", 1805 => "10101011", 1806 => "01001111", 1808 => "11110010", 1809 => "01111101", 1810 => "10010100", 1811 => "01011001", 1812 => "11110011", 1813 => "00111110", 1814 => "00010010", 1817 => "01111101", 1819 => "01011001", 1820 => "11100010", 1821 => "01011010", 1822 => "11010110", 1823 => "01111111", 1824 => "01111000", 1825 => "10010001", 1827 => "10001001", 1829 => "10010010", 1831 => "10000110", 1832 => "11000011", 1835 => "11001011", 1837 => "11001001", 1838 => "00101001", 1839 => "01000110", 1840 => "11011111", 1842 => "11001100", 1843 => "11100010", 1844 => "10111111", 1845 => "11100111", 1846 => "01011100", 1847 => "00000100", 1848 => "00010100", 1849 => "11100000", 1851 => "11001000", 1853 => "01101011", 1855 => "00100110", 1856 => "00000011", 1857 => "00101101", 1858 => "00001110", 1860 => "11001101", 1861 => "01111101", 1862 => "00010001", 1864 => "11110000", 1867 => "00011011", 1868 => "00100101", 1869 => "00000100", 1870 => "01101011", 1872 => "00001011", 1873 => "10011100", 1874 => "01101001", 1875 => "10011001", 1876 => "11011000", 1877 => "00111000", 1878 => "01101101", 1880 => "00110101", 1881 => "10111001", 1882 => "11000001", 1884 => "01111101", 1886 => "10000111", 1887 => "10111111", 1888 => "01001001", 1889 => "01010110", 1891 => "01010011", 1892 => "11100001", 1893 => "11010111", 1894 => "10010100", 1895 => "10110001", 1898 => "01011011", 1899 => "10110001", 1901 => "11100011", 1902 => "01000011", 1903 => "11111010", 1904 => "00000010", 1906 => "01110001", 1907 => "01111011", 1908 => "01100011", 1910 => "00100000", 1912 => "00001010", 1913 => "01001010", 1914 => "01101011", 1915 => "01110011", 1916 => "00000010", 1917 => "10110001", 1918 => "11110010", 1920 => "10011111", 1922 => "00000011", 1925 => "10000101", 1927 => "01010001", 1928 => "01100101", 1929 => "01001110", 1930 => "11110101", 1931 => "00010000", 1932 => "01110101", 1933 => "01010001", 1934 => "11100010", 1935 => "00001101", 1936 => "11010001", 1937 => "01011000", 1938 => "00011100", 1939 => "00101011", 1941 => "11011000", 1942 => "01111011", 1943 => "11010111", 1944 => "01101001", 1945 => "00011111", 1946 => "01100101", 1947 => "10101101", 1949 => "10101001", 1950 => "10000000", 1951 => "11011111", 1953 => "10111111", 1954 => "10000011", 1956 => "00010100", 1957 => "01110100", 1958 => "10010000", 1959 => "11100010", 1962 => "00100001", 1963 => "11011101", 1964 => "10011111", 1965 => "11000011", 1966 => "10000101", 1967 => "10010101", 1968 => "00000101", 1969 => "00101011", 1973 => "00100111", 1974 => "11001010", 1980 => "11101110", 1981 => "01001001", 1983 => "00011111", 1986 => "00110000", 1988 => "11111010", 1989 => "00001111", 1990 => "01000101", 1991 => "11100001", 1992 => "11001110", 1996 => "11110011", 1998 => "00010001", 2000 => "10111010", 2001 => "01110000", 2002 => "11010111", 2004 => "01110011", 2005 => "11011010", 2006 => "01010010", 2008 => "01011111", 2010 => "11100000", 2011 => "01100101", 2012 => "00011010", 2014 => "00111100", 2016 => "01010010", 2017 => "11100000", 2018 => "11001011", 2019 => "11100101", 2021 => "11101110", 2023 => "01100010", 2024 => "00111101", 2025 => "10000101", 2026 => "01111000", 2027 => "00101101", 2029 => "11001010", 2030 => "00111100", 2031 => "11000101", 2032 => "11110111", 2033 => "01101101", 2034 => "01000111", 2035 => "10011001", 2037 => "11011110", 2038 => "01111101", 2040 => "11000011", 2041 => "10101101", 2042 => "11110001", 2044 => "10011100", 2045 => "01001101", 2046 => "11111101", 2048 => "10010000", 2049 => "01010011", 2050 => "00010010", 2051 => "00111000", 2052 => "01110000", 2053 => "01010111", 2055 => "11011001", 2058 => "00011011", 2060 => "10001110", 2061 => "11100001", 2062 => "00000101", 2065 => "00101010", 2066 => "01101101", 2067 => "10100100", 2068 => "10010011", 2070 => "11010011", 2071 => "01111011", 2072 => "10111010", 2073 => "11010001", 2075 => "10111001", 2076 => "01110011", 2077 => "10011110", 2078 => "10001101", 2079 => "01110001", 2081 => "01101110", 2082 => "01000010", 2084 => "00100100", 2085 => "11110011", 2086 => "11101111", 2087 => "11101100", 2088 => "11111000", 2089 => "00000010", 2090 => "01010100", 2091 => "01100110", 2093 => "00101010", 2094 => "00100100", 2095 => "10100011", 2096 => "11100111", 2097 => "01000101", 2098 => "01110000", 2100 => "00101111", 2101 => "01000101", 2103 => "11011101", 2104 => "01011000", 2106 => "10101011", 2107 => "01001010", 2109 => "01001010", 2110 => "01001110", 2112 => "01000100", 2113 => "11111111", 2114 => "10100001", 2115 => "10101100", 2116 => "00111111", 2117 => "10110100", 2118 => "10010101", 2119 => "11000011", 2120 => "11110001", 2121 => "11111110", 2122 => "00010100", 2124 => "00010100", 2125 => "01000010", 2126 => "00101000", 2128 => "10100111", 2129 => "10001100", 2131 => "01101010", 2132 => "01001101", 2135 => "01100111", 2136 => "01001111", 2140 => "11010110", 2141 => "10110111", 2142 => "11111001", 2143 => "00100001", 2144 => "00001100", 2145 => "01111001", 2146 => "10101011", 2149 => "10100010", 2150 => "01100001", 2152 => "11000011", 2153 => "01010101", 2154 => "01011111", 2155 => "10010011", 2156 => "00110011", 2158 => "01101001", 2160 => "00001000", 2162 => "00011001", 2163 => "10101001", 2165 => "10110000", 2166 => "11100001", 2167 => "00111001", 2169 => "11000011", 2170 => "10000111", 2171 => "00111101", 2172 => "00001100", 2175 => "00011100", 2176 => "00000111", 2177 => "11101101", 2178 => "10100011", 2179 => "10100101", 2180 => "01000010", 2181 => "01110001", 2182 => "01011100", 2183 => "10010101", 2184 => "11010111", 2185 => "11100110", 2189 => "11011111", 2190 => "11111101", 2191 => "11010110", 2192 => "00101011", 2193 => "11000001", 2194 => "11010010", 2195 => "11100001", 2196 => "10000100", 2199 => "11110010", 2200 => "01011010", 2201 => "01100010", 2204 => "01010001", 2205 => "11110101", 2206 => "01000100", 2208 => "10111011", 2209 => "10111010", 2210 => "11101111", 2212 => "11100001", 2214 => "11101101", 2215 => "01011111", 2217 => "00111110", 2218 => "00110001", 2219 => "10001100", 2220 => "00100100", 2221 => "10111111", 2222 => "00110001", 2223 => "00100110", 2224 => "10000011", 2227 => "00011111", 2229 => "00110011", 2230 => "00010111", 2233 => "10001001", 2235 => "01000100", 2236 => "11111111", 2237 => "01111110", 2239 => "10100000", 2240 => "10000110", 2242 => "11111110", 2243 => "01000010", 2244 => "11111011", 2247 => "11010001", 2248 => "01001011", 2249 => "01111111", 2250 => "00001101", 2251 => "10000110", 2252 => "11011101", 2253 => "10110111", 2254 => "11010001", 2256 => "11001111", 2257 => "11101010", 2259 => "11010111", 2261 => "00100101", 2262 => "01000111", 2263 => "10001100", 2264 => "10000010", 2265 => "00010100", 2266 => "00101111", 2267 => "01011111", 2268 => "10011101", 2270 => "00111110", 2271 => "01111001", 2273 => "01101100", 2274 => "10111101", 2275 => "00000011", 2276 => "11011101", 2277 => "11110000", 2278 => "11000000", 2279 => "11010010", 2280 => "11101010", 2282 => "01100101", 2283 => "11111100", 2284 => "00111011", 2285 => "10111010", 2286 => "01011111", 2288 => "10001010", 2290 => "11110000", 2291 => "11111101", 2292 => "00010110", 2293 => "01111110", 2294 => "10101110", 2295 => "01011011", 2296 => "11010000", 2297 => "10100100", 2298 => "11100111", 2299 => "00011001", 2302 => "00001101", 2303 => "01100101", 2304 => "10001100", 2307 => "00000101", 2308 => "01001000", 2309 => "00111100", 2312 => "01011101", 2313 => "11011000", 2315 => "10000110", 2316 => "10111011", 2317 => "01010010", 2318 => "01000010", 2320 => "01011101", 2322 => "11001010", 2324 => "10000100", 2326 => "00100111", 2328 => "10101001", 2329 => "11101111", 2331 => "00111000", 2333 => "01100001", 2334 => "01110100", 2335 => "11001000", 2337 => "11110110", 2338 => "00010110", 2339 => "11101011", 2340 => "01000001", 2342 => "01000010", 2343 => "01011001", 2345 => "01001110", 2346 => "01111010", 2347 => "11011100", 2348 => "00100100", 2349 => "10011010", 2350 => "11101111", 2351 => "00100011", 2352 => "10110011", 2353 => "01010011", 2354 => "10111011", 2355 => "10011000", 2356 => "11111010", 2359 => "01101000", 2360 => "11101001", 2361 => "11000010", 2366 => "11101100", 2370 => "01010011", 2371 => "11110101", 2373 => "01001011", 2375 => "01100010", 2376 => "10100000", 2377 => "11100010", 2378 => "11111111", 2380 => "10101011", 2383 => "00110000", 2384 => "00110011", 2385 => "01001111", 2387 => "00001010", 2388 => "01101011", 2389 => "11011011", 2390 => "10100101", 2391 => "01011100", 2393 => "11010111", 2396 => "01110100", 2397 => "10001111", 2401 => "11110100", 2402 => "11000011", 2407 => "01001010", 2408 => "01101001", 2409 => "10110011", 2410 => "01111000", 2412 => "00011010", 2413 => "10110010", 2416 => "01111010", 2417 => "10011011", 2420 => "10101111", 2421 => "00000001", 2423 => "01011011", 2424 => "10010011", 2425 => "10010100", 2429 => "01011110", 2430 => "00001110", 2431 => "00010001", 2432 => "11110010", 2433 => "10011001", 2434 => "11000000", 2435 => "00111101", 2437 => "01110000", 2438 => "00110000", 2440 => "01010000", 2441 => "11100100", 2442 => "00110100", 2443 => "11100110", 2444 => "01101011", 2445 => "01000010", 2446 => "01101100", 2448 => "00110101", 2449 => "00011011", 2450 => "10010111", 2452 => "11010111", 2453 => "00010011", 2454 => "11110100", 2455 => "10010000", 2456 => "11000011", 2457 => "11110010", 2458 => "01111000", 2460 => "10011011", 2461 => "10000000", 2462 => "10000011", 2463 => "10010110", 2466 => "01100101", 2468 => "01011101", 2469 => "10101110", 2470 => "00010100", 2471 => "00111100", 2472 => "10010011", 2473 => "00001111", 2474 => "00011010", 2476 => "00000001", 2477 => "00010110", 2479 => "01001001", 2480 => "01111000", 2481 => "10000100", 2483 => "11000111", 2484 => "10111011", 2485 => "01010000", 2487 => "00111010", 2488 => "11111001", 2489 => "10100111", 2490 => "11100001", 2492 => "11000000", 2493 => "00101001", 2494 => "11000111", 2496 => "11000111", 2497 => "00100101", 2498 => "01101101", 2499 => "00011000", 2500 => "11101101", 2501 => "11111000", 2502 => "01001101", 2504 => "10110111", 2505 => "01010110", 2507 => "01001010", 2508 => "01011100", 2509 => "01100110", 2510 => "11110110", 2512 => "10101101", 2514 => "10110000", 2515 => "00000001", 2516 => "11100000", 2517 => "10101111", 2518 => "11010001", 2519 => "10110000", 2521 => "11011111", 2522 => "10100101", 2523 => "00111101", 2524 => "11100111", 2526 => "10111001", 2529 => "11011100", 2531 => "00011000", 2532 => "00111110", 2535 => "00100101", 2538 => "10100011", 2539 => "11010001", 2540 => "00001001", 2541 => "10000101", 2542 => "11000110", 2543 => "10110001", 2544 => "00001111", 2545 => "00000010", 2547 => "00110000", 2549 => "10011001", 2550 => "01001010", 2551 => "11010011", 2552 => "10011000", 2553 => "00010001", 2555 => "00011001", 2556 => "01010000", 2557 => "01001011", 2559 => "00101100", 2560 => "11101001", 2561 => "00100000", 2562 => "10110111", 2563 => "10100010", 2564 => "11110110", 2565 => "00011101", 2566 => "11101010", 2567 => "11010111", 2569 => "00111010", 2570 => "10001001", 2571 => "00010011", 2572 => "10010111", 2573 => "00100111", 2575 => "11101010", 2576 => "00010110", 2577 => "00001010", 2579 => "10010100", 2581 => "10001101", 2582 => "01101111", 2583 => "11000001", 2584 => "11101000", 2588 => "11011011", 2589 => "10111011", 2590 => "10010101", 2591 => "00001100", 2592 => "10011010", 2594 => "11100001", 2597 => "11011100", 2598 => "11001100", 2600 => "11110101", 2601 => "10101000", 2603 => "01001110", 2604 => "00100000", 2605 => "00110000", 2606 => "11000001", 2608 => "00100100", 2609 => "11110011", 2610 => "01001010", 2611 => "01111011", 2613 => "11000101", 2614 => "11100000", 2615 => "00000010", 2616 => "11101001", 2618 => "10000000", 2619 => "11111010", 2620 => "10010111", 2621 => "11101110", 2622 => "01100100", 2623 => "10101001", 2625 => "11001110", 2629 => "11010000", 2630 => "10011111", 2631 => "10011001", 2632 => "00101000", 2633 => "01100011", 2634 => "11111101", 2635 => "00000101", 2636 => "00000010", 2637 => "10101101", 2638 => "00000010", 2639 => "01110001", 2640 => "00010111", 2642 => "00010011", 2643 => "11101011", 2644 => "10011010", 2646 => "11111011", 2647 => "11100000", 2648 => "10010111", 2649 => "11110001", 2650 => "11100100", 2651 => "11011101", 2653 => "01101110", 2654 => "11110000", 2655 => "10110111", 2656 => "00100010", 2657 => "01111111", 2659 => "01100011", 2660 => "11000100", 2661 => "10010000", 2662 => "01000000", 2663 => "11001001", 2665 => "00011011", 2666 => "01011100", 2667 => "01010100", 2668 => "10100000", 2670 => "00100100", 2673 => "00101011", 2674 => "10110010", 2676 => "11011000", 2677 => "01010111", 2678 => "00011011", 2679 => "11010001", 2680 => "10001101", 2681 => "00111101", 2683 => "00010101", 2685 => "10000100", 2686 => "10001111", 2687 => "10011111", 2688 => "10111001", 2691 => "00100000", 2693 => "00101111", 2694 => "11110110", 2696 => "00011011", 2697 => "00111111", 2698 => "11111111", 2699 => "01001111", 2700 => "11010000", 2701 => "11010100", 2702 => "11100101", 2704 => "10001011", 2705 => "01110001", 2706 => "00101111", 2707 => "10010011", 2708 => "11000011", 2709 => "11000011", 2710 => "11010001", 2711 => "10010111", 2712 => "11010011", 2715 => "10111010", 2717 => "10111101", 2718 => "10001011", 2719 => "00101011", 2720 => "10000010", 2724 => "00000100", 2726 => "10001000", 2727 => "01011011", 2728 => "11010011", 2729 => "00111101", 2730 => "01000110", 2731 => "11110100", 2732 => "11110110", 2733 => "10011100", 2735 => "00011001", 2736 => "01110011", 2737 => "01111010", 2738 => "00010110", 2739 => "01011001", 2741 => "10011001", 2743 => "10011101", 2744 => "01011001", 2746 => "10101100", 2747 => "11011010", 2749 => "01101000", 2751 => "00110011", 2753 => "11111110", 2754 => "10001101", 2757 => "00100010", 2758 => "11001110", 2759 => "00000010", 2760 => "11100000", 2761 => "01000000", 2762 => "00000011", 2763 => "01010001", 2764 => "00100001", 2767 => "00010000", 2768 => "10000000", 2769 => "10001000", 2774 => "10111000", 2776 => "11101000", 2777 => "10010101", 2778 => "10101101", 2779 => "01110011", 2781 => "11001100", 2782 => "00011100", 2783 => "11011110", 2784 => "10011111", 2785 => "11110101", 2786 => "01001001", 2787 => "10110010", 2788 => "10101010", 2789 => "11001111", 2790 => "10001100", 2791 => "10101010", 2792 => "10111100", 2793 => "10010110", 2795 => "00100011", 2796 => "11001111", 2797 => "00010000", 2798 => "01101001", 2799 => "10000010", 2801 => "00010010", 2803 => "01010011", 2805 => "01011100", 2806 => "10011001", 2807 => "11000100", 2808 => "00011000", 2810 => "11110111", 2812 => "01101000", 2814 => "01011000", 2815 => "11101010", 2817 => "10110000", 2818 => "10111101", 2819 => "11111100", 2821 => "00101110", 2822 => "01111111", 2823 => "11011111", 2824 => "11010100", 2825 => "10001101", 2826 => "10000100", 2827 => "00000111", 2828 => "01001110", 2829 => "00010110", 2830 => "00010011", 2831 => "01111110", 2836 => "00010100", 2839 => "11010010", 2840 => "11010100", 2842 => "00010000", 2844 => "01001010", 2845 => "11000111", 2846 => "10000111", 2847 => "11010000", 2848 => "00001101", 2849 => "01000011", 2850 => "01010000", 2851 => "00011010", 2852 => "10011001", 2853 => "00111011", 2854 => "11001111", 2856 => "00100001", 2858 => "00110101", 2859 => "10110000", 2860 => "00010110", 2863 => "11000101", 2867 => "00110111", 2868 => "10001010", 2869 => "11101010", 2870 => "11100101", 2871 => "00011101", 2872 => "01010000", 2873 => "01100010", 2874 => "10000010", 2876 => "11101101", 2878 => "11100110", 2879 => "00100010", 2881 => "11100111", 2882 => "00101000", 2883 => "11011000", 2884 => "10101000", 2885 => "11110100", 2886 => "01001010", 2888 => "00101011", 2889 => "01011011", 2891 => "00010111", 2893 => "10011110", 2894 => "01010000", 2896 => "01000111", 2897 => "10100101", 2898 => "00001000", 2899 => "01011110", 2901 => "00100101", 2903 => "10001101", 2904 => "10111001", 2905 => "11111110", 2907 => "11110011", 2908 => "10000000", 2909 => "11101010", 2910 => "10001111", 2911 => "00110101", 2912 => "11111101", 2913 => "01111000", 2914 => "00010010", 2915 => "01010001", 2916 => "00101001", 2917 => "00001111", 2918 => "10010110", 2919 => "00000010", 2921 => "11101010", 2923 => "11101010", 2924 => "01110010", 2925 => "01110100", 2927 => "00101110", 2928 => "11001101", 2929 => "01001110", 2931 => "00001111", 2932 => "10001011", 2933 => "11010101", 2934 => "10111110", 2935 => "11001000", 2936 => "01010010", 2939 => "00100110", 2940 => "10101101", 2941 => "00001010", 2942 => "11100111", 2944 => "00000110", 2945 => "01000111", 2946 => "11000110", 2947 => "00011011", 2948 => "01110011", 2950 => "00111010", 2951 => "00010110", 2952 => "10100011", 2954 => "11010001", 2957 => "00110100", 2958 => "11101101", 2959 => "01110010", 2961 => "00001000", 2962 => "01010111", 2963 => "01000001", 2966 => "10000001", 2969 => "00110010", 2970 => "01111001", 2971 => "10100110", 2973 => "00110001", 2976 => "10110010", 2977 => "10101110", 2978 => "00000010", 2979 => "10000001", 2981 => "00100000", 2982 => "01010011", 2983 => "11110101", 2985 => "01010101", 2986 => "00110000", 2987 => "10100001", 2988 => "00011101", 2989 => "01010111", 2990 => "11010101", 2992 => "11100010", 2994 => "11100111", 2995 => "00001100", 2996 => "10001010", 2997 => "00011100", 2999 => "01111110", 3002 => "11101010", 3003 => "10001100", 3004 => "00011010", 3005 => "10110011", 3007 => "10111000", 3008 => "11010011", 3009 => "01101011", 3010 => "11110000", 3011 => "00011000", 3012 => "00101001", 3013 => "11011101", 3014 => "11100101", 3015 => "10110011", 3016 => "11011001", 3018 => "10100100", 3019 => "11000110", 3020 => "00001111", 3021 => "11000110", 3022 => "00011111", 3024 => "10001111", 3025 => "11011000", 3027 => "00110101", 3028 => "01111000", 3029 => "01001000", 3031 => "01011110", 3032 => "10001001", 3033 => "01010001", 3034 => "01110010", 3035 => "10110011", 3039 => "00100000", 3040 => "10101011", 3041 => "10111110", 3042 => "01110011", 3043 => "11011010", 3044 => "01111000", 3045 => "10001010", 3046 => "01100001", 3047 => "00000010", 3048 => "01111110", 3050 => "10100101", 3052 => "10001010", 3053 => "00001010", 3054 => "00000101", 3055 => "10000110", 3057 => "11000101", 3058 => "11100110", 3059 => "10001111", 3060 => "01010110", 3061 => "01101001", 3062 => "10101100", 3063 => "10111110", 3064 => "10110001", 3066 => "10001110", 3067 => "00001111", 3068 => "11000101", 3069 => "10111001", 3071 => "01101010", 3073 => "00011100", 3074 => "01100010", 3075 => "10000011", 3076 => "11110111", 3077 => "10101000", 3078 => "10101010", 3079 => "10001000", 3080 => "01000001", 3081 => "11011011", 3082 => "10111110", 3083 => "10110000", 3085 => "11100110", 3086 => "01111010", 3087 => "10111101", 3088 => "10010111", 3089 => "00000010", 3091 => "00001100", 3095 => "10101110", 3096 => "01001010", 3097 => "11000000", 3098 => "10111001", 3100 => "10111011", 3103 => "11011000", 3105 => "11111011", 3106 => "11101001", 3107 => "11100111", 3108 => "01101010", 3110 => "10011010", 3111 => "00111010", 3112 => "00011101", 3113 => "00001100", 3114 => "11000100", 3115 => "10001101", 3116 => "11011001", 3117 => "10101101", 3118 => "10001010", 3120 => "00101101", 3121 => "10111010", 3122 => "11000010", 3124 => "10001100", 3125 => "01110110", 3126 => "11001110", 3128 => "01000001", 3130 => "01110010", 3131 => "00110000", 3132 => "11100000", 3133 => "00010101", 3134 => "10101010", 3135 => "00111110", 3137 => "10010000", 3138 => "01100101", 3139 => "00001000", 3141 => "11101100", 3142 => "00111111", 3144 => "11010110", 3145 => "01010111", 3146 => "01000100", 3147 => "00001110", 3148 => "00101100", 3149 => "01011100", 3150 => "00010100", 3151 => "11000010", 3152 => "11001110", 3153 => "00100100", 3156 => "10111100", 3158 => "00111111", 3159 => "10111110", 3160 => "11000101", 3162 => "10010110", 3163 => "00011111", 3164 => "10011011", 3165 => "00010100", 3166 => "11110110", 3168 => "11101110", 3169 => "11010010", 3170 => "11001111", 3173 => "10110100", 3174 => "01011010", 3176 => "01100111", 3178 => "11110100", 3179 => "10110010", 3180 => "11110010", 3181 => "00000100", 3182 => "01100011", 3184 => "01010101", 3186 => "11000000", 3187 => "01110001", 3188 => "11110000", 3189 => "11111101", 3190 => "11001001", 3191 => "11100011", 3192 => "00100001", 3194 => "01011110", 3195 => "01011010", 3196 => "10101010", 3197 => "11000101", 3198 => "10001001", 3199 => "00000100", 3200 => "00010110", 3202 => "11111011", 3203 => "01111001", 3204 => "01110010", 3207 => "01101111", 3208 => "10110000", 3209 => "01011011", 3210 => "11011001", 3211 => "11011001", 3212 => "11010000", 3213 => "10100010", 3214 => "11111110", 3215 => "01011110", 3218 => "10110011", 3219 => "11011011", 3220 => "00010101", 3221 => "01010110", 3222 => "10000101", 3223 => "00101000", 3224 => "10011010", 3226 => "01011100", 3227 => "10001100", 3228 => "10000101", 3229 => "00101101", 3230 => "00000001", 3231 => "11111101", 3232 => "10011001", 3235 => "10011000", 3236 => "01000100", 3237 => "00111010", 3238 => "11110010", 3240 => "11000101", 3241 => "00101011", 3243 => "00011011", 3245 => "01100111", 3247 => "01011100", 3248 => "10011111", 3249 => "11001011", 3250 => "00000110", 3251 => "11000100", 3252 => "00000001", 3253 => "10011110", 3255 => "00010011", 3256 => "11100011", 3257 => "11100010", 3258 => "00011001", 3259 => "00000111", 3260 => "00110001", 3261 => "10101111", 3262 => "11100000", 3263 => "11001101", 3264 => "00010001", 3265 => "11000110", 3266 => "01111001", 3267 => "11010010", 3269 => "11100110", 3271 => "11000110", 3272 => "01100000", 3273 => "00010010", 3276 => "10011011", 3277 => "11000100", 3278 => "01110001", 3279 => "10010000", 3280 => "01000010", 3282 => "11001111", 3283 => "11010100", 3284 => "10001101", 3287 => "01011110", 3289 => "01110011", 3290 => "11100110", 3291 => "11100010", 3293 => "11101111", 3294 => "10001011", 3295 => "00101111", 3296 => "10110111", 3298 => "11001001", 3299 => "10100101", 3304 => "00010000", 3305 => "01110000", 3307 => "00100110", 3308 => "01010000", 3310 => "00010001", 3311 => "11100101", 3312 => "10010010", 3313 => "10000101", 3315 => "11100001", 3318 => "01010011", 3319 => "00001010", 3320 => "11010100", 3324 => "01101110", 3326 => "01111100", 3327 => "11110010", 3328 => "11010111", 3329 => "01111110", 3330 => "10101101", 3333 => "11000011", 3334 => "11011101", 3335 => "00111001", 3336 => "10000110", 3337 => "11001110", 3338 => "01101110", 3340 => "10000011", 3341 => "10000111", 3342 => "10111101", 3343 => "00111110", 3344 => "00110010", 3345 => "01000000", 3346 => "10011001", 3347 => "01110000", 3348 => "11001101", 3349 => "01101100", 3351 => "00110001", 3352 => "10010000", 3353 => "10001011", 3354 => "11100001", 3355 => "00101110", 3356 => "01111011", 3357 => "11110100", 3358 => "00000010", 3360 => "00010010", 3361 => "01101110", 3362 => "11010010", 3364 => "11000100", 3366 => "00010011", 3367 => "11010010", 3368 => "11101101", 3369 => "11001000", 3370 => "00100000", 3371 => "00101001", 3372 => "00011001", 3373 => "11001010", 3374 => "10001100", 3378 => "10010100", 3379 => "10100010", 3380 => "00011111", 3381 => "00101111", 3382 => "10010011", 3383 => "00011000", 3384 => "01011101", 3387 => "00011010", 3388 => "00000001", 3389 => "01000010", 3391 => "10101011", 3392 => "10001000", 3393 => "00100001", 3394 => "10001100", 3395 => "00100110", 3396 => "00000110", 3398 => "01111000", 3399 => "11101110", 3401 => "00011010", 3402 => "10000101", 3406 => "11111000", 3407 => "10011010", 3411 => "01100101", 3412 => "00010110", 3415 => "00000111", 3416 => "11000000", 3417 => "11010010", 3419 => "00101000", 3421 => "01101101", 3423 => "00101101", 3424 => "11100100", 3425 => "01010100", 3426 => "00010010", 3427 => "10101111", 3429 => "11010111", 3430 => "00000110", 3431 => "11000011", 3432 => "00001101", 3433 => "00100100", 3434 => "11001100", 3436 => "01011101", 3437 => "01111011", 3438 => "10010000", 3440 => "11101100", 3441 => "11010110", 3442 => "01011011", 3443 => "11011010", 3444 => "11101010", 3445 => "11110011", 3446 => "01110001", 3447 => "00011011", 3448 => "01001011", 3449 => "01011101", 3450 => "10000010", 3451 => "10001010", 3452 => "10000110", 3453 => "11110000", 3455 => "00110000", 3456 => "11001110", 3457 => "10011010", 3458 => "10101101", 3459 => "11001001", 3460 => "00010011", 3461 => "01100010", 3462 => "11110111", 3463 => "01110011", 3464 => "00000001", 3465 => "10011101", 3466 => "10100111", 3467 => "10110001", 3468 => "11011111", 3469 => "01110010", 3470 => "11101110", 3471 => "11000111", 3472 => "11010010", 3473 => "11111010", 3475 => "00100011", 3476 => "00001110", 3478 => "00111010", 3479 => "11110100", 3482 => "10011000", 3484 => "01110101", 3485 => "01001011", 3486 => "01110000", 3488 => "10100011", 3489 => "10011011", 3491 => "11001111", 3494 => "10110010", 3498 => "10001000", 3499 => "01100110", 3500 => "01011111", 3502 => "11000001", 3504 => "11111011", 3506 => "01011110", 3507 => "10011111", 3508 => "00011001", 3510 => "10000011", 3511 => "11100010", 3512 => "01010010", 3513 => "10001011", 3515 => "01100110", 3517 => "10100101", 3519 => "00000001", 3520 => "10011101", 3521 => "01011000", 3522 => "11100010", 3526 => "10100001", 3527 => "00100110", 3531 => "00111111", 3532 => "00111011", 3533 => "10010001", 3536 => "00100001", 3537 => "10100101", 3538 => "10001111", 3539 => "10011010", 3541 => "10001100", 3543 => "11101100", 3544 => "00011101", 3547 => "10110001", 3548 => "00101001", 3550 => "10001000", 3551 => "01011001", 3552 => "10011110", 3554 => "10000010", 3555 => "01010111", 3557 => "10011001", 3558 => "10100001", 3559 => "11010011", 3561 => "11011000", 3568 => "00111001", 3569 => "01010110", 3571 => "01011110", 3572 => "11011010", 3573 => "00100101", 3577 => "11110011", 3579 => "10001101", 3586 => "00110011", 3587 => "01111100", 3590 => "01110110", 3591 => "11000101", 3593 => "10110111", 3594 => "00111011", 3595 => "01010111", 3597 => "01111001", 3601 => "01101110", 3602 => "00010110", 3603 => "11011110", 3605 => "11110000", 3611 => "00111111", 3612 => "10100110", 3613 => "01000000", 3614 => "10110100", 3616 => "00010111", 3618 => "01011110", 3620 => "11000101", 3622 => "11100000", 3624 => "10010100", 3625 => "10010000", 3627 => "10101101", 3628 => "11101100", 3634 => "00100101", 3637 => "00111000", 3639 => "01101001", 3640 => "11010100", 3641 => "10000010", 3644 => "00010100", 3648 => "00111111", 3649 => "10111110", 3653 => "01111101", 3657 => "00100111", 3658 => "10011001", 3660 => "10101001", 3662 => "00111011", 3663 => "01101000", 3665 => "11011101", 3666 => "00101111", 3667 => "01000001", 3669 => "10010011", 3670 => "01011101", 3673 => "11010111", 3677 => "01110001", 3680 => "01011101", 3681 => "10111101", 3685 => "01011100", 3687 => "10111100", 3688 => "01101001", 3689 => "01100110", 3691 => "11101110", 3698 => "01011010", 3699 => "00111101", 3701 => "01100100", 3702 => "11000111", 3705 => "11011101", 3707 => "00000001", 3712 => "00010110", 3713 => "01011111", 3714 => "00101100", 3718 => "00110110", 3723 => "11101010", 3726 => "00010010", 3727 => "00010010", 3729 => "10011111", 3731 => "01111010", 3732 => "00001111", 3735 => "01111010", 3737 => "00011111", 3740 => "01001010", 3744 => "00010000", 3746 => "10111111", 3747 => "00011111", 3748 => "01011000", 3751 => "00011001", 3753 => "01001000", 3759 => "00011101", 3760 => "01110100", 3762 => "10010011", 3763 => "00100010", 3768 => "10000011", 3769 => "01101110", 3770 => "01010101", 3772 => "10001011", 3773 => "00000111", 3774 => "10111011", 3775 => "00011101", 3777 => "01011110", 3778 => "10011101", 3779 => "11001101", 3780 => "10110100", 3781 => "11101101", 3782 => "01100011", 3784 => "00111100", 3786 => "00001101", 3787 => "10100010", 3788 => "10000011", 3789 => "00101101", 3791 => "10110000", 3792 => "01100000", 3793 => "01110100", 3794 => "10000000", 3796 => "10010110", 3797 => "11011111", 3798 => "11110100", 3800 => "00110101", 3803 => "01001100", 3804 => "10111101", 3807 => "01011001", 3809 => "01100111", 3812 => "00001011", 3814 => "11101110", 3818 => "10010100", 3819 => "00011011", 3820 => "01001011", 3821 => "10000011", 3824 => "10010101", 3825 => "10101000", 3826 => "01101011", 3828 => "10110000", 3835 => "01010100", 3839 => "01110011", 3840 => "10001001", 3842 => "11000011", 3843 => "01110110", 3844 => "01001101", 3845 => "10000011", 3847 => "10110011", 3853 => "10010010", 3854 => "11000111", 3857 => "11001101", 3861 => "11001010", 3864 => "00010001", 3866 => "10000010", 3867 => "10110100", 3869 => "10010010", 3870 => "01101011", 3872 => "00101110", 3873 => "10100110", 3874 => "00011001", 3875 => "00001011", 3876 => "11000011", 3879 => "10001011", 3881 => "11010000", 3883 => "11110000", 3884 => "11010000", 3885 => "10010001", 3887 => "11110011", 3888 => "10000101", 3893 => "00001010", 3894 => "00110010", 3895 => "10101011", 3897 => "11011101", 3898 => "00110101", 3904 => "00001100", 3905 => "00000101", 3906 => "11000111", 3907 => "10110010", 3913 => "10010011", 3914 => "01101000", 3917 => "00011010", 3918 => "01101111", 3921 => "01011110", 3922 => "11111000", 3923 => "01011011", 3924 => "00010100", 3927 => "11010110", 3928 => "11010101", 3931 => "10101001", 3932 => "01010111", 3933 => "00001101", 3937 => "11010000", 3938 => "10100110", 3939 => "11110110", 3940 => "10100011", 3941 => "11111101", 3947 => "11011101", 3950 => "11001001", 3952 => "01010100", 3956 => "10011100", 3957 => "11101001", 3958 => "10111001", 3962 => "01110101", 3963 => "01110110", 3964 => "10111101", 3965 => "10001110", 3966 => "11010011", 3967 => "00100100", 3971 => "10000110", 3972 => "01001100", 3973 => "11111001", 3975 => "11111011", 3977 => "00101101", 3978 => "00110111", 3981 => "00100001", 3982 => "01010011", 3983 => "10100010", 3984 => "11000110", 3987 => "11101100", 3988 => "11011001", 3990 => "10110101", 3991 => "00011101", 3995 => "10100001", 3996 => "10000101", 4006 => "00101011", 4008 => "01001000", 4011 => "00011010", 4012 => "00111111", 4013 => "01001001", 4016 => "01110000", 4017 => "10111001", 4020 => "11000001", 4023 => "00011011", 4024 => "10110100", 4025 => "11001001", 4026 => "10001011", 4029 => "11010111", 4032 => "11000110", 4040 => "11010110", 4043 => "11010100", 4046 => "11001110", 4048 => "11110111", 4049 => "10001000", 4053 => "00110000", 4055 => "01011010", 4056 => "01101011", 4058 => "11101000", 4060 => "01011010", 4061 => "00100010", 4062 => "11010111", 4063 => "11010100", 4064 => "01101101", 4067 => "11110000", 4068 => "01010000", 4071 => "01011011", 4073 => "00110010", 4074 => "10111010", 4075 => "00100001", 4076 => "00011111", 4082 => "00000111", 4083 => "10101100", 4084 => "01001111", 4086 => "01110000", 4090 => "10010111", 4092 => "11000011", 4093 => "10001000", 4094 => "10100100", 4096 => "01011001", 4098 => "01101101", 4101 => "01111010", 4106 => "11101110", 4108 => "11010001", 4110 => "10000010", 4112 => "11111000", 4114 => "01101110", 4115 => "10101111", 4118 => "00111011", 4120 => "00100000", 4121 => "01000011", 4122 => "01111110", 4123 => "00010101", 4126 => "00001111", 4131 => "11101101", 4134 => "11011000", 4135 => "00010111", 4136 => "10110111", 4141 => "10110000", 4143 => "11101100", 4144 => "00000011", 4149 => "11001101", 4151 => "01111100", 4152 => "11001101", 4154 => "10100101", 4155 => "00101111", 4156 => "10111001", 4157 => "10110011", 4158 => "00101110", 4160 => "11001001", 4163 => "11100001", 4164 => "00100000", 4165 => "11010101", 4166 => "01011100", 4169 => "01001110", 4173 => "01100100", 4175 => "11001000", 4176 => "10110010", 4178 => "01001000", 4181 => "01100100", 4182 => "00101010", 4184 => "11011100", 4189 => "00100100", 4193 => "10100100", 4194 => "01111100", 4195 => "11101001", 4196 => "10101100", 4200 => "01100110", 4201 => "01010010", 4202 => "10011101", 4205 => "01000110", 4207 => "11010001", 4212 => "01001001", 4214 => "01010010", 4216 => "01011111", 4218 => "01100111", 4219 => "10100110", 4220 => "10111101", 4223 => "10101110", 4224 => "10111111", 4226 => "11011011", 4227 => "11001011", 4231 => "10000010", 4232 => "01010101", 4236 => "11111100", 4238 => "01100100", 4239 => "10010011", 4242 => "11001011", 4251 => "01100101", 4253 => "00111001", 4255 => "01111011", 4259 => "10000001", 4260 => "10111100", 4261 => "01000110", 4264 => "11011000", 4265 => "00011010", 4266 => "01001011", 4267 => "01111100", 4268 => "01010001", 4269 => "10011101", 4271 => "10100001", 4276 => "01011011", 4277 => "11110000", 4282 => "10001110", 4284 => "11001100", 4288 => "11001111", 4291 => "01011010", 4293 => "11000000", 4294 => "00101100", 4297 => "11100100", 4298 => "10010011", 4300 => "11100001", 4301 => "10101111", 4304 => "01100110", 4305 => "11100111", 4307 => "11011111", 4308 => "00110101", 4311 => "11001110", 4312 => "10111000", 4314 => "10000000", 4315 => "01111100", 4316 => "01010111", 4318 => "10111110", 4320 => "01110000", 4321 => "01000000", 4323 => "10110100", 4331 => "11000110", 4332 => "00011000", 4334 => "11010001", 4336 => "10000110", 4337 => "00000101", 4338 => "11000111", 4341 => "11111001", 4343 => "00111111", 4346 => "11101100", 4347 => "01111110", 4348 => "11101110", 4351 => "11001011", 4360 => "11101110", 4364 => "11110011", 4365 => "11111001", 4368 => "01110010", 4372 => "00001000", 4373 => "01010011", 4375 => "00100100", 4377 => "01111100", 4381 => "11000001", 4385 => "00011101", 4386 => "11010101", 4388 => "01100000", 4389 => "10011000", 4390 => "00101101", 4392 => "01001001", 4396 => "01001110", 4397 => "11011011", 4402 => "01010000", 4405 => "11110111", 4406 => "00100000", 4408 => "00011000", 4409 => "11111000", 4411 => "00110000", 4414 => "11001100", 4415 => "01100101", 4416 => "01010010", 4420 => "10000111", 4421 => "10100011", 4422 => "11101100", 4423 => "00010000", 4424 => "01001100", 4426 => "00011100", 4428 => "00001001", 4429 => "00001011", 4431 => "00000100", 4432 => "11100111", 4434 => "11010100", 4435 => "11111110", 4437 => "10001110", 4445 => "11011011", 4448 => "10101110", 4449 => "00010110", 4450 => "10100011", 4452 => "11101100", 4453 => "00011110", 4454 => "10011011", 4457 => "00101001", 4458 => "00010000", 4459 => "11111011", 4462 => "10101110", 4466 => "01110100", 4467 => "10000100", 4468 => "11110110", 4470 => "00111010", 4473 => "01011001", 4474 => "11100001", 4478 => "11101100", 4479 => "10001010", 4482 => "01011000", 4485 => "10011100", 4488 => "01001110", 4490 => "11110001", 4492 => "01110100", 4493 => "10010010", 4494 => "00111101", 4499 => "11100010", 4500 => "10011000", 4503 => "01101111", 4504 => "10111000", 4506 => "01011110", 4507 => "11100111", 4509 => "10010110", 4510 => "00100100", 4513 => "00000100", 4517 => "01100111", 4522 => "01101011", 4523 => "10101100", 4526 => "11001000", 4532 => "10000011", 4533 => "00010010", 4534 => "00001111", 4538 => "11110101", 4540 => "10001111", 4542 => "11000010", 4543 => "11111001", 4544 => "11011101", 4546 => "01100010", 4547 => "10111100", 4548 => "00110010", 4550 => "11001010", 4552 => "10000110", 4554 => "10111001", 4555 => "11100000", 4556 => "11111010", 4559 => "10010110", 4560 => "10010011", 4562 => "00010100", 4563 => "11000010", 4564 => "00010101", 4566 => "01101111", 4568 => "00001010", 4570 => "01001110", 4571 => "10011001", 4574 => "00101000", 4576 => "11000000", 4577 => "00000001", 4578 => "01000011", 4580 => "10001101", 4582 => "00011101", 4583 => "11001110", 4584 => "11011111", 4585 => "00110100", 4589 => "00100010", 4594 => "11111011", 4596 => "10101101", 4597 => "10001110", 4598 => "00001010", 4599 => "10101000", 4603 => "00111011", 4604 => "11000011", 4605 => "00101110", 4606 => "11011100", 4607 => "10011001", 4609 => "01100011", 4610 => "11011001", 4611 => "10101111", 4612 => "11110011", 4613 => "00110001", 4614 => "10101011", 4616 => "11010100", 4622 => "00001100", 4623 => "10101010", 4624 => "11111000", 4628 => "01111110", 4630 => "10000100", 4631 => "01010000", 4633 => "10000101", 4634 => "01001001", 4637 => "01011111", 4639 => "11111110", 4640 => "11110000", 4642 => "11011100", 4644 => "11101001", 4648 => "10011110", 4651 => "01000001", 4652 => "10001011", 4653 => "11111110", 4655 => "11110001", 4656 => "01011010", 4659 => "01100100", 4660 => "11100011", 4666 => "01010111", 4668 => "01100010", 4672 => "11110011", 4673 => "11000111", 4674 => "11000100", 4676 => "11110001", 4679 => "11010001", 4682 => "00100110", 4683 => "00100001", 4685 => "11100100", 4686 => "10110111", 4687 => "11000010", 4689 => "10011110", 4691 => "01001000", 4692 => "10000101", 4694 => "10010001", 4695 => "01000101", 4699 => "01001110", 4700 => "00011110", 4702 => "11101100", 4707 => "10001011", 4709 => "10011101", 4710 => "11010110", 4711 => "10011011", 4714 => "01101010", 4716 => "10111111", 4717 => "11101011", 4719 => "01000100", 4720 => "01010111", 4721 => "00110100", 4722 => "10101110", 4727 => "00101101", 4731 => "11101101", 4735 => "00100110", 4737 => "11010111", 4741 => "10110010", 4742 => "10001000", 4743 => "01000010", 4747 => "01001101", 4748 => "10101100", 4749 => "01011000", 4750 => "00111001", 4753 => "10101001", 4754 => "10101100", 4756 => "00100001", 4758 => "01001010", 4761 => "01010011", 4762 => "10011011", 4767 => "01101010", 4769 => "11001100", 4771 => "00011011", 4774 => "01001110", 4777 => "00110010", 4779 => "10011011", 4780 => "00011001", 4783 => "11111100", 4786 => "10100000", 4787 => "01000111", 4788 => "00001101", 4795 => "10011101", 4797 => "00111010", 4798 => "01001100", 4800 => "01010000", 4801 => "01000111", 4802 => "00110101", 4803 => "00101101", 4806 => "10110011", 4808 => "00111000", 4810 => "11000010", 4812 => "01001110", 4814 => "00111100", 4815 => "10100110", 4817 => "10010110", 4821 => "11010100", 4823 => "10010101", 4824 => "00110111", 4826 => "01100101", 4827 => "00111110", 4831 => "11101001", 4833 => "10111101", 4834 => "10101101", 4835 => "00010001", 4836 => "01101011", 4838 => "11100101", 4841 => "11000010", 4843 => "10000100", 4844 => "10100000", 4845 => "00101111", 4847 => "01101100", 4849 => "00101010", 4851 => "01110011", 4856 => "01000000", 4857 => "00111110", 4859 => "10011100", 4862 => "01001000", 4864 => "00110011", 4867 => "11100000", 4868 => "01011011", 4870 => "11101010", 4873 => "10000101", 4874 => "11010101", 4877 => "10100100", 4878 => "11001010", 4881 => "11111110", 4882 => "10011011", 4883 => "10100001", 4887 => "11010101", 4888 => "01000010", 4889 => "11000110", 4893 => "01110010", 4894 => "01011100", 4896 => "11000000", 4899 => "10100001", 4907 => "11000000", 4910 => "00000100", 4917 => "00001000", 4918 => "10000101", 4920 => "00010101", 4921 => "11010010", 4922 => "10100010", 4926 => "01000100", 4927 => "11110000", 4930 => "10000001", 4932 => "10010100", 4935 => "01110110", 4936 => "11001101", 4937 => "01110011", 4939 => "11111110", 4940 => "10110111", 4941 => "11101101", 4945 => "10000011", 4948 => "01010110", 4949 => "00001010", 4954 => "00000100", 4956 => "00010111", 4961 => "00001110", 4962 => "00110100", 4963 => "00110011", 4966 => "01111100", 4967 => "10100000", 4968 => "01000011", 4975 => "01100100", 4977 => "11100001", 4982 => "11000000", 4983 => "00100100", 4984 => "01110110", 4986 => "11110101", 4989 => "01110101", 4991 => "11011110", 4995 => "11100011", 4997 => "10111010", 4998 => "00111011", 4999 => "10110100", 5000 => "01011001", 5002 => "11010100", 5003 => "01011000", 5005 => "11100011", 5007 => "01101100", 5008 => "00101011", 5013 => "01011100", 5018 => "10101001", 5020 => "10011111", 5021 => "00000111", 5024 => "00011010", 5025 => "10101011", 5026 => "00001010", 5029 => "11111001", 5031 => "00100110", 5033 => "01001100", 5034 => "00111010", 5035 => "10001110", 5038 => "10011100", 5040 => "11110111", 5042 => "11000111", 5043 => "01101110", 5045 => "01010000", 5047 => "01100100", 5053 => "01011011", 5054 => "11100001", 5055 => "00100001", 5062 => "00100100", 5064 => "00111110", 5065 => "00101101", 5067 => "01010111", 5069 => "01001100", 5071 => "01000100", 5073 => "00101110", 5075 => "00110100", 5076 => "10011010", 5077 => "10100111", 5078 => "01100111", 5079 => "00001001", 5080 => "11011100", 5082 => "00100111", 5083 => "11000001", 5084 => "01110110", 5085 => "00110110", 5086 => "01101010", 5096 => "01111110", 5100 => "00010100", 5101 => "01001000", 5102 => "11111011", 5103 => "10110011", 5104 => "01101000", 5105 => "10100000", 5106 => "10101011", 5108 => "00111001", 5110 => "11000010", 5111 => "01100100", 5112 => "00111011", 5113 => "10010011", 5114 => "10110100", 5115 => "11000111", 5116 => "11000101", 5117 => "10011111", 5120 => "01100111", 5121 => "10001100", 5122 => "11110100", 5126 => "01111001", 5128 => "01111001", 5130 => "01100011", 5135 => "00011000", 5136 => "11000011", 5137 => "01110100", 5139 => "10001000", 5140 => "01111011", 5142 => "11100100", 5145 => "11110001", 5147 => "00100000", 5149 => "11001100", 5150 => "11011011", 5152 => "01111010", 5153 => "10100000", 5154 => "11010011", 5155 => "00001011", 5158 => "00100101", 5159 => "11111000", 5162 => "10001000", 5164 => "11011111", 5165 => "00111010", 5168 => "00011010", 5170 => "10010111", 5171 => "00110101", 5172 => "10110101", 5174 => "11001111", 5175 => "11001001", 5176 => "10011110", 5178 => "00110010", 5179 => "11010100", 5180 => "11001110", 5181 => "11011101", 5184 => "10000100", 5185 => "01100010", 5187 => "01101001", 5188 => "01111010", 5190 => "11110101", 5191 => "01011001", 5192 => "10101000", 5196 => "00010001", 5197 => "01110111", 5201 => "00010110", 5202 => "01010110", 5206 => "00000110", 5207 => "00111100", 5208 => "01010110", 5209 => "00100100", 5213 => "11001111", 5215 => "00100011", 5216 => "10101011", 5221 => "11100001", 5225 => "00110000", 5226 => "01101010", 5227 => "10011010", 5233 => "10111011", 5235 => "00101100", 5237 => "11000010", 5238 => "11111001", 5239 => "01011101", 5242 => "00110011", 5245 => "11001010", 5246 => "11010000", 5249 => "11111110", 5250 => "11100011", 5253 => "10100011", 5254 => "10001111", 5256 => "01100000", 5257 => "01001010", 5263 => "10010101", 5266 => "11110000", 5267 => "10101001", 5270 => "10111011", 5272 => "11100001", 5273 => "00101000", 5275 => "00111100", 5285 => "01101111", 5286 => "01110110", 5290 => "01010011", 5291 => "01000100", 5293 => "01010000", 5296 => "01111001", 5297 => "00100001", 5303 => "01111000", 5306 => "01110110", 5307 => "01010101", 5308 => "11110101", 5310 => "01111010", 5313 => "11111001", 5321 => "00011001", 5323 => "01111011", 5324 => "11011001", 5328 => "11011011", 5330 => "00001001", 5333 => "10110001", 5336 => "01010001", 5337 => "01110011", 5339 => "11100011", 5340 => "11001010", 5341 => "10111000", 5343 => "01001101", 5344 => "00110101", 5345 => "11001111", 5346 => "10000010", 5347 => "01010101", 5348 => "00111101", 5350 => "10100100", 5355 => "10100111", 5356 => "10010001", 5357 => "10010011", 5359 => "10111100", 5360 => "00100011", 5362 => "11001111", 5365 => "01111001", 5366 => "00001000", 5368 => "11011110", 5369 => "00110100", 5370 => "00000101", 5372 => "01011001", 5373 => "00011100", 5374 => "01111010", 5376 => "10000101", 5380 => "01110000", 5381 => "01101100", 5382 => "10110010", 5384 => "11110111", 5385 => "00111101", 5388 => "10000011", 5389 => "10011110", 5390 => "10111011", 5395 => "10010111", 5398 => "00011100", 5401 => "00000010", 5402 => "10000101", 5405 => "10010111", 5406 => "11101110", 5407 => "10010110", 5408 => "00101110", 5411 => "00011111", 5413 => "11001000", 5414 => "00111001", 5415 => "01011010", 5419 => "01010000", 5420 => "10000100", 5421 => "00011011", 5423 => "11110011", 5426 => "11000000", 5427 => "00001100", 5428 => "00111110", 5430 => "01101100", 5431 => "01011000", 5433 => "00011100", 5435 => "00110110", 5436 => "00011001", 5437 => "11001000", 5438 => "10001000", 5440 => "10110010", 5443 => "11111111", 5444 => "11101100", 5446 => "11001111", 5447 => "01111001", 5448 => "11000111", 5451 => "10101001", 5455 => "11011111", 5456 => "01110001", 5459 => "11010010", 5460 => "01010110", 5464 => "11001110", 5465 => "01001110", 5466 => "10111001", 5467 => "11101001", 5469 => "00100000", 5470 => "10111110", 5472 => "00101100", 5473 => "01011110", 5476 => "01010111", 5477 => "11000010", 5480 => "10010000", 5482 => "11101110", 5484 => "10111011", 5486 => "10010110", 5492 => "01111001", 5493 => "10001110", 5494 => "00000010", 5497 => "11010100", 5500 => "00101111", 5502 => "11001001", 5503 => "10010101", 5507 => "00100100", 5509 => "00000100", 5511 => "01000100", 5513 => "11111111", 5514 => "10010001", 5516 => "01111101", 5518 => "11110010", 5519 => "00001010", 5520 => "11011010", 5524 => "10000000", 5525 => "11000010", 5526 => "11111000", 5527 => "10110100", 5533 => "00010010", 5537 => "11101101", 5538 => "00011010", 5539 => "11001011", 5540 => "10101011", 5541 => "11111011", 5542 => "01010111", 5544 => "10000111", 5545 => "10000011", 5546 => "00011100", 5549 => "10110011", 5551 => "11101010", 5557 => "11000100", 5558 => "00101111", 5559 => "11100111", 5560 => "10100000", 5561 => "10000100", 5562 => "10001101", 5565 => "11011100", 5567 => "10011110", 5570 => "01010111", 5571 => "11011001", 5572 => "01010110", 5573 => "10111110", 5575 => "11000010", 5576 => "10110101", 5577 => "01010100", 5578 => "01011010", 5582 => "11010010", 5584 => "10011100", 5586 => "11010000", 5589 => "11000111", 5590 => "10001101", 5591 => "10011101", 5592 => "10011100", 5594 => "01000010", 5595 => "11000101", 5597 => "11010011", 5599 => "01011110", 5603 => "01100010", 5605 => "01110100", 5606 => "11011000", 5607 => "11001001", 5609 => "01011001", 5611 => "01100011", 5612 => "00011100", 5614 => "10000101", 5615 => "01110010", 5620 => "01110000", 5621 => "01001010", 5623 => "11011001", 5627 => "10011111", 5630 => "01010111", 5631 => "11100111", 5633 => "01010111", 5639 => "10111011", 5640 => "11001011", 5641 => "01100101", 5643 => "00101010", 5645 => "00011000", 5646 => "11110011", 5648 => "00011111", 5649 => "10000011", 5651 => "10001010", 5653 => "01011101", 5654 => "11100001", 5656 => "00011111", 5657 => "10010101", 5658 => "01010010", 5659 => "11111000", 5660 => "00111010", 5662 => "01100100", 5664 => "11101010", 5665 => "01111011", 5667 => "11000001", 5668 => "01101100", 5669 => "11100110", 5670 => "00111010", 5671 => "00011011", 5675 => "00100000", 5676 => "11100001", 5677 => "00110011", 5681 => "01001010", 5683 => "00010101", 5684 => "00000010", 5687 => "00011111", 5688 => "00111001", 5689 => "10000110", 5690 => "10001010", 5692 => "10011001", 5694 => "01011011", 5697 => "11001110", 5698 => "11000000", 5705 => "01000011", 5706 => "00011100", 5710 => "00000011", 5714 => "00000001", 5717 => "00110100", 5719 => "11000011", 5720 => "11110100", 5722 => "01101101", 5724 => "00010100", 5728 => "10100001", 5729 => "01000000", 5730 => "10000000", 5734 => "00010110", 5736 => "01110110", 5737 => "00001100", 5744 => "11000100", 5745 => "11011110", 5746 => "00001111", 5747 => "01101101", 5749 => "11011001", 5752 => "10010110", 5754 => "10111000", 5755 => "10101110", 5756 => "00101001", 5762 => "00000100", 5763 => "11011111", 5767 => "00011111", 5768 => "11101011", 5771 => "01011110", 5772 => "01100000", 5773 => "10111001", 5778 => "00111001", 5779 => "10110110", 5783 => "11001110", 5784 => "01101111", 5785 => "10000110", 5791 => "00110110", 5792 => "01111010", 5793 => "00011111", 5794 => "11010001", 5795 => "10001010", 5800 => "01010010", 5809 => "10011100", 5811 => "11010110", 5813 => "01111100", 5814 => "10100000", 5820 => "00100010", 5821 => "11101100", 5822 => "11011000", 5826 => "01101000", 5827 => "11000011", 5829 => "01100000", 5830 => "11110001", 5831 => "00111111", 5835 => "10000010", 5837 => "00011100", 5840 => "11100010", 5841 => "11100001", 5842 => "11001011", 5844 => "00001100", 5845 => "11101011", 5848 => "10111101", 5849 => "10000100", 5852 => "10010100", 5854 => "00011001", 5855 => "11100101", 5857 => "01000000", 5859 => "00001010", 5862 => "10110001", 5866 => "00010010", 5868 => "11001001", 5871 => "10000111", 5881 => "11011100", 5884 => "01010011", 5885 => "11110011", 5889 => "01101010", 5893 => "01110010", 5897 => "11011101", 5898 => "00001011", 5899 => "11101011", 5900 => "11000010", 5902 => "01101011", 5906 => "10110110", 5907 => "00111011", 5908 => "00001101", 5909 => "00111011", 5911 => "11100001", 5912 => "11110110", 5914 => "11010111", 5917 => "10000011", 5918 => "01011001", 5920 => "11000111", 5923 => "00011001", 5924 => "01010010", 5927 => "10001011", 5928 => "00100111", 5929 => "11100010", 5932 => "01101101", 5935 => "10100001", 5936 => "00101111", 5937 => "11100001", 5940 => "01101011", 5941 => "01110111", 5943 => "01111011", 5944 => "01101010", 5945 => "01101101", 5948 => "00010011", 5950 => "10110011", 5952 => "01011110", 5955 => "10010101", 5957 => "00101100", 5959 => "01110111", 5961 => "10101010", 5962 => "00010001", 5963 => "10100011", 5965 => "00110011", 5966 => "11010001", 5974 => "10001100", 5976 => "10010110", 5977 => "10111010", 5978 => "11011011", 5980 => "10100111", 5982 => "00011000", 5987 => "10101011", 5989 => "00101110", 5990 => "11001110", 5992 => "11011101", 5995 => "10100011", 5996 => "01000110", 5997 => "11111010", 5998 => "00010001", 6000 => "00111111", 6002 => "01000111", 6003 => "00101001", 6007 => "11100011", 6008 => "11001010", 6009 => "00001000", 6010 => "00010000", 6011 => "10000111", 6014 => "01111010", 6015 => "10101100", 6016 => "00111100", 6017 => "11011010", 6020 => "10100100", 6022 => "01011000", 6025 => "01101101", 6026 => "10010100", 6029 => "00001111", 6030 => "11010000", 6031 => "01111100", 6032 => "01011111", 6037 => "00000111", 6039 => "00010001", 6040 => "11010101", 6041 => "00100101", 6044 => "00010100", 6045 => "01000100", 6047 => "00110101", 6048 => "01100111", 6052 => "01111111", 6055 => "10101110", 6056 => "00010101", 6059 => "01101111", 6060 => "10001001", 6061 => "10110111", 6062 => "00101011", 6063 => "11111000", 6065 => "01011100", 6066 => "00011000", 6068 => "00010011", 6069 => "01101000", 6073 => "01010001", 6075 => "01100110", 6076 => "11100111", 6077 => "10111101", 6078 => "00010101", 6079 => "10111011", 6083 => "11101010", 6085 => "11000011", 6087 => "00100011", 6088 => "10001011", 6091 => "10000001", 6093 => "11010110", 6095 => "11010001", 6096 => "00100001", 6097 => "01110011", 6098 => "01000110", 6101 => "10000111", 6104 => "00010100", 6106 => "00010000", 6107 => "11010100", 6110 => "01001100", 6112 => "11101101", 6113 => "01100100", 6119 => "10110100", 6122 => "00000111", 6123 => "10110001", 6127 => "00110101", 6128 => "00101011", 6130 => "10001101", 6131 => "00000001", 6132 => "11010101", 6138 => "10011000", 6139 => "01100110", 6142 => "01110101", 6145 => "11010111", 6146 => "00010101", 6147 => "10000000", 6151 => "10101001", 6153 => "00110110", 6155 => "00000001", 6157 => "00111110", 6159 => "00101010", 6162 => "10100001", 6163 => "00110101", 6164 => "10011111", 6166 => "10001100", 6167 => "01110000", 6168 => "00100001", 6169 => "00111111", 6175 => "10000111", 6176 => "11100100", 6178 => "10010011", 6180 => "01110111", 6183 => "10100010", 6184 => "00111000", 6185 => "10011010", 6187 => "01101110", 6188 => "11100100", 6190 => "10010111", 6191 => "10111011", 6192 => "11001101", 6196 => "11110111", 6197 => "01000101", 6198 => "10101110", 6199 => "11011101", 6200 => "00110101", 6201 => "01111110", 6203 => "11100001", 6205 => "10100101", 6207 => "01001101", 6208 => "01110100", 6211 => "00110010", 6212 => "10010100", 6213 => "01001010", 6214 => "00100011", 6215 => "00010100", 6218 => "00000101", 6219 => "10011001", 6221 => "11001101", 6222 => "00000011", 6223 => "11001010", 6226 => "11010011", 6227 => "00110101", 6228 => "00101101", 6229 => "01000001", 6233 => "00000001", 6236 => "11000011", 6238 => "00001001", 6241 => "01011101", 6242 => "01110100", 6249 => "10101001", 6254 => "11001010", 6256 => "01010000", 6257 => "00001000", 6259 => "11101001", 6260 => "10100110", 6261 => "00010001", 6263 => "01100001", 6264 => "10111101", 6265 => "11001011", 6266 => "11011000", 6269 => "01101000", 6271 => "10001100", 6276 => "10010010", 6277 => "11000100", 6280 => "01111110", 6281 => "11100011", 6282 => "10100001", 6283 => "01111011", 6284 => "11101010", 6287 => "01001110", 6290 => "00011000", 6296 => "11011010", 6298 => "10011101", 6299 => "11101000", 6303 => "11101101", 6306 => "11110001", 6308 => "00100100", 6310 => "01011001", 6314 => "11001100", 6315 => "10110010", 6317 => "01101101", 6325 => "11010001", 6326 => "10000110", 6327 => "10000111", 6330 => "00000110", 6331 => "00110110", 6336 => "10101100", 6340 => "11111101", 6343 => "00100000", 6344 => "11010100", 6345 => "11000001", 6347 => "01011000", 6351 => "00001001", 6352 => "10110011", 6353 => "11100101", 6355 => "10011101", 6356 => "00000011", 6357 => "11101111", 6358 => "01111111", 6359 => "00001010", 6362 => "11101011", 6363 => "00101011", 6367 => "11000011", 6368 => "11110000", 6370 => "01100101", 6372 => "10100000", 6376 => "11100101", 6377 => "10010110", 6380 => "10010101", 6382 => "01100101", 6383 => "00011001", 6384 => "01011001", 6386 => "10110111", 6389 => "10000111", 6390 => "00000101", 6391 => "11101110", 6393 => "01001000", 6396 => "00011010", 6400 => "01001100", 6401 => "10000000", 6405 => "10000101", 6406 => "11110000", 6407 => "01010010", 6408 => "01111100", 6410 => "11011100", 6412 => "10001011", 6413 => "10010011", 6415 => "11010011", 6416 => "01111101", 6419 => "11001101", 6420 => "01101000", 6421 => "01011110", 6424 => "10100110", 6425 => "01111001", 6429 => "01001111", 6431 => "10010011", 6432 => "00000111", 6436 => "00111101", 6437 => "11111111", 6438 => "01000010", 6439 => "10101001", 6441 => "10100001", 6442 => "01111110", 6448 => "11110110", 6449 => "11111101", 6450 => "00100100", 6451 => "01010110", 6455 => "01111001", 6461 => "01010011", 6462 => "00001111", 6463 => "11100100", 6465 => "00011100", 6466 => "00100110", 6467 => "11000011", 6468 => "01010000", 6469 => "00111010", 6472 => "01110100", 6474 => "00010011", 6476 => "10010011", 6477 => "00100010", 6479 => "10011111", 6483 => "11010100", 6488 => "11011010", 6490 => "11011101", 6491 => "01100000", 6492 => "11001010", 6493 => "01000001", 6494 => "10000000", 6497 => "11010011", 6499 => "00110000", 6500 => "10110010", 6503 => "00011000", 6507 => "11011100", 6508 => "11100011", 6509 => "10000100", 6512 => "11001100", 6515 => "11010011", 6520 => "01101101", 6522 => "00111101", 6524 => "10100110", 6525 => "11110011", 6529 => "00100001", 6533 => "10111010", 6536 => "01000011", 6538 => "10001100", 6539 => "01100010", 6541 => "11100010", 6542 => "01110101", 6544 => "11010001", 6548 => "11111111", 6550 => "01110000", 6551 => "01100111", 6553 => "00010110", 6555 => "01010011", 6556 => "11001011", 6558 => "10000000", 6560 => "01010101", 6561 => "11100101", 6562 => "01100010", 6564 => "11000111", 6565 => "00011101", 6566 => "10101000", 6570 => "10001011", 6572 => "01111111", 6573 => "00100110", 6576 => "11100100", 6578 => "00010111", 6583 => "01100001", 6585 => "01101111", 6586 => "01110110", 6588 => "10000001", 6589 => "10001001", 6591 => "10111101", 6595 => "11100010", 6597 => "01011110", 6598 => "11111101", 6602 => "10101010", 6606 => "10101000", 6608 => "10011110", 6611 => "00101000", 6612 => "00110101", 6614 => "10010100", 6615 => "01100111", 6619 => "01101100", 6623 => "00101100", 6624 => "10100100", 6625 => "11010001", 6631 => "01111000", 6632 => "10001010", 6633 => "10110010", 6634 => "10001011", 6635 => "11000101", 6638 => "11000000", 6640 => "01110111", 6643 => "11010110", 6644 => "01101110", 6645 => "10011101", 6649 => "00000101", 6651 => "01101110", 6653 => "10100000", 6654 => "00001100", 6655 => "01001000", 6656 => "01000000", 6657 => "01000100", 6660 => "10111001", 6661 => "10100000", 6662 => "00011100", 6665 => "10010100", 6667 => "10100010", 6668 => "00010101", 6669 => "10110111", 6675 => "11010010", 6677 => "10011011", 6680 => "00100101", 6682 => "01010011", 6683 => "10011001", 6684 => "00111010", 6686 => "00000001", 6687 => "10001101", 6688 => "00011100", 6690 => "01111111", 6691 => "10000000", 6692 => "10011000", 6694 => "11010100", 6695 => "10000110", 6704 => "00000110", 6705 => "10110110", 6706 => "01100010", 6709 => "00000111", 6714 => "11001111", 6715 => "00001000", 6716 => "11110100", 6718 => "01100010", 6719 => "01000000", 6720 => "10111111", 6721 => "11100101", 6722 => "11001101", 6725 => "10111011", 6728 => "01100100", 6731 => "11110001", 6732 => "11011011", 6734 => "10111000", 6735 => "01000001", 6739 => "11011000", 6740 => "00010101", 6741 => "10011110", 6746 => "01011101", 6747 => "01011001", 6748 => "00000101", 6750 => "01001111", 6754 => "10101011", 6756 => "00100000", 6764 => "00011001", 6765 => "11101001", 6768 => "01100011", 6769 => "10000010", 6770 => "11001011", 6772 => "11111111", 6773 => "01100100", 6775 => "00011010", 6778 => "11000010", 6779 => "10110111", 6781 => "00010001", 6782 => "10111111", 6784 => "00100100", 6785 => "00001101", 6788 => "00101100", 6793 => "10111010", 6796 => "11001000", 6797 => "01100111", 6798 => "11001111", 6803 => "00100011", 6804 => "10100101", 6805 => "11001010", 6806 => "00100111", 6809 => "10100011", 6810 => "01010110", 6811 => "11010010", 6815 => "01010100", 6816 => "11101001", 6817 => "01010000", 6818 => "11000001", 6822 => "00000101", 6823 => "00111101", 6827 => "10100010", 6828 => "10100010", 6830 => "10100111", 6833 => "01110101", 6838 => "11100001", 6840 => "01110100", 6843 => "10000001", 6849 => "11010110", 6850 => "00001000", 6851 => "01111100", 6852 => "11001111", 6854 => "11100100", 6856 => "01110011", 6857 => "10111101", 6858 => "01011100", 6860 => "00001011", 6861 => "00011110", 6863 => "00111100", 6867 => "00010100", 6874 => "00101100", 6875 => "01000011", 6876 => "11111001", 6877 => "01101110", 6879 => "01000011", 6882 => "00111000", 6887 => "00111011", 6888 => "11000110", 6890 => "00001101", 6892 => "01111000", 6898 => "01000010", 6901 => "10010001", 6904 => "00010101", 6905 => "10111101", 6909 => "00111110", 6911 => "10110001", 6914 => "01100110", 6916 => "00001100", 6917 => "00000101", 6918 => "10010000", 6919 => "01010110", 6921 => "00010100", 6922 => "11001000", 6923 => "00111100", 6924 => "10000010", 6926 => "00111100", 6928 => "10010110", 6931 => "11011011", 6933 => "01010111", 6936 => "01110110", 6938 => "01110011", 6939 => "01011001", 6940 => "00111100", 6941 => "11111101", 6945 => "01001110", 6946 => "10111000", 6947 => "00100100", 6952 => "11010011", 6954 => "11001010", 6957 => "10101100", 6962 => "10010000", 6963 => "01011100", 6964 => "11011111", 6965 => "01000000", 6966 => "01101111", 6968 => "00100100", 6969 => "01101010", 6970 => "11100110", 6974 => "01110110", 6975 => "00001000", 6977 => "11111010", 6980 => "01001110", 6984 => "10001111", 6985 => "11001111", 6986 => "01101011", 6987 => "11000011", 6988 => "11001011", 6989 => "11101001", 6990 => "00110001", 6994 => "11000011", 6996 => "00110011", 6997 => "00000110", 6999 => "10110101", 7000 => "11101110", 7001 => "01101001", 7004 => "10010101", 7007 => "01000010", 7008 => "10101101", 7009 => "11111100", 7010 => "11101001", 7011 => "10000100", 7013 => "10001101", 7014 => "01111111", 7015 => "10101101", 7016 => "00110101", 7017 => "00011100", 7021 => "10010000", 7025 => "00000110", 7028 => "11010000", 7029 => "00011011", 7033 => "11000100", 7037 => "10000100", 7039 => "00010111", 7042 => "10100110", 7045 => "01010011", 7046 => "10110111", 7047 => "11110001", 7048 => "10001110", 7050 => "10000010", 7051 => "01010000", 7053 => "10010101", 7054 => "01110100", 7055 => "01111011", 7057 => "00000100", 7059 => "01000100", 7062 => "11111111", 7068 => "11111010", 7069 => "11111000", 7070 => "01111111", 7071 => "01000010", 7074 => "00000011", 7077 => "00010110", 7078 => "00110000", 7080 => "01111110", 7081 => "10000101", 7088 => "11001010", 7089 => "00011001", 7090 => "10010111", 7091 => "11110010", 7093 => "11010011", 7094 => "01011110", 7095 => "00000100", 7096 => "00001001", 7098 => "01010000", 7099 => "10000101", 7113 => "11011101", 7114 => "10100101", 7116 => "00111110", 7119 => "01100001", 7121 => "00101101", 7122 => "01100100", 7125 => "10111001", 7126 => "10110010", 7128 => "11010110", 7131 => "10101110", 7132 => "01110100", 7133 => "00011010", 7135 => "11111110", 7138 => "10010001", 7140 => "00100011", 7142 => "00100100", 7143 => "01110111", 7145 => "01000000", 7150 => "00110010", 7153 => "01000000", 7155 => "11010110", 7158 => "01100111", 7161 => "10101010", 7164 => "00100010", 7167 => "01110111", 7168 => "01111101", 7171 => "01101101", 7177 => "01110000", 7178 => "00101101", 7184 => "10110011", 7185 => "01001001", 7187 => "01100000", 7188 => "01010001", 7191 => "11110111", 7192 => "01110101", 7194 => "11100100", 7196 => "01111100", 7197 => "10111011", 7200 => "00100110", 7201 => "00101100", 7202 => "10001111", 7203 => "00110100", 7206 => "11110000", 7210 => "00101011", 7211 => "11111010", 7212 => "00101111", 7215 => "01111110", 7216 => "11001100", 7217 => "00111011", 7220 => "00010100", 7221 => "10110011", 7223 => "10011100", 7224 => "01110011", 7225 => "01011101", 7230 => "11010010", 7234 => "00100110", 7235 => "10011011", 7236 => "10000110", 7237 => "01000111", 7239 => "10111111", 7240 => "11111100", 7241 => "11111001", 7246 => "11001001", 7249 => "11001111", 7251 => "10000110", 7253 => "10001110", 7257 => "01111100", 7261 => "10111110", 7262 => "00101101", 7263 => "00001010", 7267 => "00100100", 7268 => "00100011", 7270 => "00011011", 7271 => "01011111", 7273 => "10010010", 7274 => "10101110", 7278 => "00110000", 7280 => "11100001", 7285 => "01100011", 7287 => "10011000", 7288 => "10000101", 7289 => "01110100", 7290 => "00101010", 7295 => "11001010", 7296 => "01000010", 7297 => "10100001", 7300 => "01101101", 7301 => "11101001", 7303 => "00111001", 7304 => "11001110", 7308 => "11000001", 7311 => "00100001", 7313 => "11101011", 7315 => "11101110", 7316 => "10011111", 7317 => "10000101", 7318 => "00010101", 7321 => "01011111", 7322 => "01100000", 7324 => "11111100", 7326 => "10010000", 7329 => "11001001", 7338 => "00010111", 7339 => "11101100", 7342 => "11000101", 7345 => "00110110", 7346 => "00010111", 7347 => "11111010", 7349 => "10101101", 7350 => "11011000", 7353 => "00000110", 7355 => "00110000", 7356 => "01001101", 7358 => "10010010", 7364 => "11010101", 7369 => "00101001", 7373 => "11101010", 7379 => "11101101", 7380 => "00100011", 7383 => "01111100", 7385 => "11110101", 7386 => "00010100", 7387 => "11100101", 7388 => "00101010", 7389 => "11111010", 7392 => "01010011", 7393 => "10000010", 7394 => "11101011", 7395 => "11010110", 7396 => "00011001", 7397 => "10111000", 7398 => "00110101", 7400 => "01000001", 7402 => "10110010", 7403 => "00001001", 7404 => "10010100", 7407 => "01111001", 7408 => "01010010", 7415 => "11010011", 7416 => "01011110", 7417 => "11010011", 7420 => "01111000", 7421 => "00001111", 7422 => "11111010", 7423 => "01100101", 7426 => "01001110", 7427 => "11010010", 7429 => "11000010", 7431 => "00011101", 7432 => "10101110", 7435 => "00101001", 7437 => "10001101", 7440 => "00101001", 7442 => "11000111", 7446 => "11001101", 7449 => "11101111", 7450 => "10110100", 7453 => "01011000", 7454 => "01100011", 7458 => "11111000", 7459 => "10111001", 7463 => "00010001", 7464 => "00001010", 7465 => "01111100", 7466 => "11011111", 7467 => "11010101", 7470 => "10010010", 7473 => "10101011", 7476 => "11100111", 7478 => "00100100", 7479 => "01110100", 7482 => "11000110", 7483 => "00101100", 7484 => "00110010", 7485 => "01010010", 7486 => "00110100", 7487 => "00101111", 7489 => "00101011", 7490 => "11010001", 7491 => "10111101", 7492 => "01110000", 7493 => "11000110", 7494 => "01000010", 7495 => "11110010", 7497 => "10001010", 7498 => "11110000", 7499 => "01100110", 7500 => "00110111", 7503 => "10001100", 7507 => "10100111", 7510 => "11101100", 7512 => "10111010", 7521 => "00010100", 7522 => "01100100", 7525 => "00111101", 7529 => "11011000", 7530 => "00011001", 7531 => "00101111", 7532 => "10110101", 7536 => "11111000", 7537 => "10110101", 7538 => "00101111", 7540 => "00001111", 7542 => "10110000", 7544 => "11011011", 7546 => "10110010", 7547 => "00010110", 7548 => "11110100", 7549 => "00100000", 7550 => "01000100", 7553 => "00000101", 7557 => "01011101", 7558 => "00010011", 7559 => "10111000", 7561 => "00101110", 7566 => "11111000", 7572 => "11000111", 7574 => "11001001", 7576 => "10101110", 7577 => "01111100", 7578 => "11111110", 7583 => "10110011", 7588 => "10111011", 7590 => "01111111", 7591 => "01001011", 7592 => "00001001", 7595 => "01110000", 7596 => "10000001", 7601 => "11110111", 7602 => "10011101", 7603 => "01000111", 7607 => "01101111", 7609 => "10111110", 7610 => "01011011", 7618 => "01100110", 7621 => "01110011", 7622 => "10111110", 7624 => "10110100", 7628 => "00101010", 7631 => "00010110", 7634 => "11101010", 7635 => "10111110", 7637 => "11111011", 7638 => "10010010", 7639 => "00100001", 7643 => "10000001", 7645 => "00110001", 7647 => "10000110", 7653 => "10100110", 7655 => "00111100", 7657 => "01010110", 7659 => "01100011", 7660 => "01110100", 7661 => "11111101", 7662 => "01001010", 7663 => "11000101", 7664 => "11110100", 7666 => "11001011", 7667 => "01000001", 7670 => "11010100", 7672 => "11111001", 7678 => "01110111", 7679 => "10100110", 7681 => "00001110", 7683 => "10001000", 7684 => "11011110", 7688 => "11001001", 7689 => "00000010", 7690 => "10101111", 7691 => "01111110", 7692 => "01100100", 7693 => "01001100", 7695 => "10010101", 7696 => "01011010", 7699 => "10010110", 7701 => "11110110", 7702 => "00000111", 7704 => "10000100", 7705 => "00111111", 7707 => "01100001", 7708 => "00110010", 7709 => "10010101", 7710 => "00111010", 7713 => "00111110", 7715 => "00011100", 7718 => "11010100", 7720 => "00100001", 7721 => "01011101", 7722 => "10101011", 7723 => "10001111", 7724 => "11101111", 7727 => "01010000", 7731 => "10011100", 7739 => "11011101", 7742 => "11101010", 7744 => "11111111", 7745 => "00111001", 7753 => "01001001", 7755 => "01111100", 7756 => "01101101", 7759 => "01000010", 7762 => "00001100", 7764 => "01010001", 7767 => "10110001", 7768 => "01110101", 7769 => "10110001", 7770 => "01010000", 7772 => "01001101", 7774 => "01000110", 7777 => "10110000", 7780 => "00001010", 7781 => "11001000", 7782 => "11010101", 7786 => "10100010", 7789 => "01111000", 7791 => "01100110", 7792 => "11110011", 7794 => "11101000", 7797 => "11101110", 7799 => "10001001", 7807 => "00110010", 7808 => "00000101", 7814 => "11111101", 7817 => "00010010", 7819 => "00111100", 7825 => "01101010", 7826 => "11111000", 7827 => "10100011", 7828 => "10101110", 7829 => "01001000", 7830 => "10101011", 7831 => "00111100", 7833 => "11000011", 7838 => "00011111", 7839 => "10010010", 7847 => "11000001", 7848 => "01000101", 7851 => "11101100", 7852 => "10010100", 7854 => "00011011", 7855 => "11110110", 7857 => "01110000", 7859 => "01110110", 7860 => "11011110", 7863 => "10000000", 7865 => "10100100", 7867 => "00010101", 7868 => "10111110", 7869 => "10101100", 7870 => "01111010", 7872 => "01011110", 7873 => "10111111", 7874 => "01000010", 7876 => "10101011", 7877 => "01111101", 7879 => "01010000", 7880 => "01011111", 7881 => "01000000", 7882 => "00100010", 7883 => "10111110", 7885 => "11011100", 7886 => "11110101", 7888 => "01101111", 7889 => "00111010", 7890 => "10101110", 7894 => "10010110", 7899 => "01000010", 7901 => "01011100", 7903 => "11110111", 7904 => "11101100", 7909 => "01000110", 7913 => "10011110", 7917 => "01011001", 7918 => "01111010", 7919 => "00010011", 7923 => "00010011", 7924 => "10111100", 7925 => "01001100", 7926 => "00100011", 7928 => "10001011", 7932 => "11011011", 7940 => "01101101", 7941 => "00101100", 7942 => "10111100", 7945 => "11011001", 7948 => "10101000", 7949 => "11001101", 7952 => "01100110", 7953 => "10011000", 7954 => "01110011", 7955 => "00000010", 7956 => "01011010", 7957 => "11110000", 7958 => "00110010", 7960 => "10011111", 7961 => "11101010", 7962 => "11011100", 7963 => "10010111", 7966 => "11111011", 7967 => "00100101", 7968 => "00100010", 7971 => "00101111", 7972 => "00001011", 7973 => "01100110", 7977 => "11010010", 7978 => "00001111", 7979 => "01110001", 7981 => "01101010", 7983 => "11100000", 7984 => "11110110", 7985 => "00111101", 7987 => "10001111", 7992 => "10001010", 7994 => "11010100", 7995 => "11000000", 7997 => "11100011", 8001 => "01001111", 8005 => "01011101", 8006 => "11110100", 8007 => "10110000", 8008 => "11000100", 8009 => "10011010", 8010 => "11011001", 8011 => "11100100", 8014 => "10011110", 8019 => "00001011", 8022 => "11001110", 8025 => "01100000", 8027 => "10000100", 8029 => "11110011", 8031 => "00010010", 8032 => "10011001", 8033 => "01010100", 8034 => "10010011", 8037 => "00011001", 8038 => "01110001", 8042 => "00010010", 8043 => "11111011", 8045 => "11101011", 8047 => "10010001", 8052 => "00010111", 8056 => "10110011", 8060 => "11010000", 8062 => "01111110", 8063 => "11110011", 8066 => "01110001", 8072 => "11001011", 8073 => "01111010", 8075 => "10010001", 8076 => "01001111", 8078 => "01010010", 8079 => "01100010", 8080 => "11001111", 8082 => "00100010", 8083 => "01010110", 8088 => "00111100", 8089 => "10111111", 8098 => "01000001", 8099 => "01001111", 8100 => "00110100", 8101 => "11000100", 8103 => "11110101", 8105 => "00101000", 8107 => "11110000", 8111 => "01101010", 8116 => "01001010", 8118 => "01000000", 8121 => "01000110", 8122 => "10010001", 8127 => "00101001", 8129 => "00100010", 8136 => "11111100", 8137 => "10011100", 8138 => "00001000", 8139 => "01110000", 8142 => "00100111", 8143 => "10110011", 8144 => "11011000", 8145 => "10011101", 8146 => "01110101", 8151 => "10110010", 8154 => "00010011", 8157 => "01011111", 8158 => "10101000", 8159 => "10011001", 8160 => "10110101", 8161 => "11110100", 8163 => "01111001", 8165 => "01010010", 8168 => "01011111", 8169 => "01111111", 8170 => "00011010", 8172 => "10111111", 8173 => "01101010", 8175 => "10110101", 8176 => "01111111", 8177 => "11011110", 8178 => "01101001", 8180 => "11001111", 8187 => "00000010", 8188 => "10000000", 8189 => "11100111", 8190 => "01110101", 8194 => "11001111", 8196 => "00101101", 8198 => "00010100", 8200 => "01101011", 8204 => "11111101", 8205 => "11000100", 8208 => "10101010", 8209 => "11101101", 8210 => "00011110", 8211 => "01110011", 8212 => "11011111", 8216 => "10000011", 8222 => "11111111", 8223 => "10000110", 8226 => "10110101", 8228 => "11010101", 8230 => "00101011", 8231 => "10011100", 8234 => "00001001", 8235 => "01110100", 8237 => "11100010", 8238 => "00010011", 8239 => "01100001", 8240 => "11000110", 8241 => "00101111", 8243 => "10001000", 8246 => "00001010", 8249 => "00011001", 8250 => "11111101", 8251 => "10001100", 8252 => "11110010", 8253 => "00100011", 8256 => "10111100", 8258 => "10001011", 8259 => "11000001", 8263 => "10110001", 8264 => "11001101", 8265 => "11010000", 8266 => "01000101", 8269 => "10101110", 8271 => "10110100", 8273 => "10010001", 8276 => "00010000", 8277 => "01101101", 8278 => "11011100", 8282 => "11000010", 8283 => "11101110", 8284 => "01111000", 8287 => "01011010", 8288 => "11101110", 8291 => "11111011", 8292 => "01110010", 8293 => "00000010", 8296 => "00101011", 8298 => "10001100", 8299 => "01001110", 8300 => "11011101", 8301 => "01100110", 8303 => "10011001", 8304 => "00000010", 8306 => "11101110", 8307 => "01101100", 8309 => "01100101", 8311 => "11010010", 8312 => "10111001", 8313 => "10001110", 8315 => "01101111", 8317 => "00111111", 8319 => "11011111", 8320 => "11110110", 8321 => "00001111", 8322 => "11101011", 8325 => "10001101", 8327 => "01011101", 8328 => "00010100", 8329 => "01101111", 8330 => "10101111", 8331 => "01000011", 8332 => "00001001", 8338 => "00110010", 8341 => "00110001", 8343 => "01011000", 8344 => "00110001", 8345 => "10000101", 8347 => "00011001", 8349 => "00101101", 8353 => "10110110", 8354 => "00000010", 8356 => "00110000", 8357 => "01010000", 8358 => "10110101", 8361 => "00011101", 8362 => "00101110", 8364 => "01000010", 8365 => "11100010", 8366 => "11010111", 8369 => "01110101", 8370 => "01001010", 8372 => "01011000", 8375 => "10111011", 8377 => "10011101", 8380 => "01001110", 8382 => "01001100", 8383 => "01110111", 8385 => "01011110", 8389 => "11110111", 8392 => "10101001", 8393 => "11011011", 8394 => "10111011", 8395 => "00011000", 8397 => "01110110", 8398 => "01001100", 8400 => "11001111", 8402 => "01110100", 8403 => "01110101", 8405 => "00011000", 8406 => "01011010", 8409 => "11111100", 8411 => "11110001", 8412 => "11101001", 8413 => "00100001", 8415 => "00111110", 8418 => "01011100", 8419 => "00101110", 8420 => "11001010", 8424 => "10001000", 8425 => "01011100", 8426 => "10101100", 8427 => "10000110", 8428 => "01111011", 8430 => "01101101", 8434 => "11110100", 8440 => "00111101", 8441 => "00111010", 8442 => "10010110", 8443 => "00011110", 8444 => "10010010", 8445 => "00100100", 8446 => "10010111", 8447 => "00100111", 8448 => "00111100", 8451 => "10111111", 8452 => "00100011", 8458 => "00010111", 8464 => "00000111", 8465 => "01001011", 8469 => "10001001", 8472 => "10011110", 8474 => "10000100", 8475 => "10100100", 8476 => "01111101", 8477 => "00100001", 8478 => "00111000", 8479 => "10001000", 8480 => "11011101", 8481 => "11101010", 8483 => "10000110", 8487 => "01011111", 8490 => "00000101", 8491 => "11110100", 8492 => "01010101", 8493 => "11101110", 8494 => "11111111", 8496 => "01000000", 8497 => "10001010", 8498 => "11100011", 8499 => "11011001", 8500 => "00001010", 8501 => "10101101", 8504 => "10001011", 8505 => "00100000", 8506 => "00000101", 8507 => "00101100", 8508 => "10111011", 8513 => "01000001", 8517 => "01001000", 8519 => "11011000", 8521 => "00011101", 8525 => "11111011", 8526 => "11001110", 8527 => "10010001", 8533 => "10111001", 8535 => "11001101", 8539 => "11011010", 8540 => "01110110", 8541 => "11110010", 8545 => "00010000", 8546 => "10100001", 8547 => "10111000", 8548 => "00000110", 8550 => "01010100", 8552 => "00110100", 8559 => "11010100", 8562 => "00100010", 8563 => "01110100", 8564 => "01100100", 8567 => "00111011", 8568 => "11001111", 8569 => "01010001", 8572 => "00101111", 8573 => "01101001", 8577 => "11000000", 8579 => "10000100", 8580 => "11010000", 8581 => "11110001", 8584 => "01000100", 8589 => "11011011", 8590 => "11101110", 8591 => "11100101", 8593 => "01000111", 8594 => "10011000", 8597 => "11101001", 8598 => "01101000", 8600 => "11010111", 8601 => "11011010", 8602 => "10101000", 8604 => "00011001", 8605 => "11000110", 8607 => "10110011", 8611 => "10101101", 8612 => "11010111", 8616 => "10110101", 8619 => "11100001", 8622 => "10110011", 8624 => "10110111", 8625 => "01111001", 8627 => "00000011", 8628 => "01100111", 8629 => "00110100", 8630 => "00101100", 8631 => "00110001", 8632 => "00101011", 8633 => "00010101", 8635 => "11100001", 8636 => "10110000", 8637 => "10001000", 8638 => "01110000", 8642 => "00111111", 8644 => "00100101", 8645 => "10000000", 8649 => "00100111", 8650 => "10100101", 8652 => "11010010", 8653 => "11111110", 8654 => "01111100", 8656 => "10001101", 8657 => "01011000", 8659 => "00001001", 8660 => "11010110", 8661 => "10011101", 8662 => "10111011", 8663 => "01111110", 8664 => "01101101", 8665 => "00110010", 8668 => "10110100", 8669 => "00100111", 8670 => "10100001", 8672 => "00100010", 8673 => "10111111", 8674 => "11001100", 8676 => "10001100", 8679 => "01110101", 8680 => "00100011", 8681 => "00010101", 8682 => "11010010", 8683 => "10011101", 8685 => "01010111", 8687 => "01100110", 8691 => "01110111", 8692 => "00000001", 8695 => "01101100", 8696 => "10001111", 8697 => "11011110", 8698 => "11011000", 8700 => "10101001", 8702 => "11010001", 8703 => "00101011", 8706 => "10101011", 8707 => "11110000", 8709 => "10100010", 8710 => "01100101", 8712 => "11111000", 8714 => "01101000", 8715 => "01000010", 8717 => "10111111", 8720 => "10010111", 8722 => "11100000", 8723 => "11001111", 8727 => "00001000", 8730 => "00000011", 8733 => "00100000", 8736 => "01001000", 8738 => "00110111", 8740 => "00001000", 8741 => "00111000", 8742 => "01111000", 8744 => "00101101", 8751 => "10011011", 8754 => "00100010", 8756 => "00011111", 8758 => "00010011", 8762 => "11000110", 8765 => "00001101", 8767 => "00111110", 8771 => "00111111", 8772 => "00110100", 8775 => "10101001", 8776 => "00110010", 8777 => "10011011", 8780 => "11011111", 8782 => "11100000", 8785 => "11001101", 8787 => "01101100", 8788 => "10011000", 8789 => "01111011", 8790 => "11100100", 8793 => "10011010", 8794 => "01100000", 8802 => "01110100", 8803 => "01010101", 8804 => "00111101", 8806 => "11111001", 8810 => "10000100", 8816 => "10000100", 8818 => "00000111", 8819 => "01001011", 8820 => "11010111", 8822 => "01111000", 8823 => "00101010", 8826 => "11101000", 8827 => "11100100", 8830 => "10110000", 8831 => "01111111", 8834 => "10100010", 8835 => "01100111", 8837 => "10000110", 8838 => "01110111", 8846 => "01000000", 8855 => "00001000", 8856 => "10111110", 8858 => "01110111", 8859 => "11000001", 8860 => "10011110", 8862 => "10111001", 8863 => "11111011", 8864 => "10001111", 8865 => "11010001", 8866 => "00111100", 8868 => "11101111", 8871 => "01010000", 8873 => "11111011", 8874 => "11001111", 8878 => "10001101", 8879 => "10000011", 8882 => "10000111", 8884 => "11010101", 8886 => "10100010", 8888 => "10110010", 8889 => "00001110", 8894 => "10100110", 8895 => "01010000", 8899 => "11100101", 8900 => "11000100", 8902 => "11100111", 8904 => "11100011", 8909 => "00010110", 8912 => "10010111", 8913 => "01010000", 8916 => "10100100", 8917 => "00011111", 8918 => "01100010", 8922 => "00101000", 8925 => "11000001", 8929 => "00010101", 8930 => "00101110", 8932 => "11010011", 8934 => "11001110", 8935 => "11110110", 8945 => "01000010", 8946 => "11000110", 8947 => "11000011", 8950 => "11001111", 8953 => "11111111", 8956 => "11101110", 8958 => "00111110", 8959 => "10011011", 8960 => "00010011", 8961 => "00110010", 8963 => "11111000", 8967 => "11001101", 8973 => "10100010", 8974 => "00110111", 8976 => "11011111", 8981 => "11011110", 8984 => "01001100", 8988 => "01011011", 8989 => "01010000", 8990 => "00100011", 8995 => "10110111", 8999 => "01011111", 9001 => "11110111", 9002 => "10101111", 9003 => "11010001", 9004 => "01000000", 9007 => "01011100", 9011 => "11100111", 9016 => "00110100", 9020 => "01000010", 9021 => "01101110", 9023 => "11100100", 9029 => "11110011", 9030 => "01001110", 9033 => "10100000", 9034 => "11000101", 9038 => "01100011", 9040 => "00110001", 9043 => "10010110", 9050 => "00000100", 9052 => "11000010", 9053 => "10001101", 9054 => "10000110", 9059 => "10110111", 9061 => "00101010", 9062 => "01101000", 9064 => "11111101", 9065 => "11010000", 9066 => "00001110", 9074 => "10111010", 9075 => "00111001", 9077 => "01011010", 9079 => "10101100", 9081 => "01110100", 9085 => "00000110", 9088 => "01000110", 9089 => "11011010", 9092 => "10110011", 9095 => "10001001", 9096 => "10111100", 9100 => "01101010", 9101 => "11101101", 9106 => "10111010", 9110 => "00111010", 9113 => "10100001", 9114 => "10001010", 9118 => "00111111", 9119 => "10111110", 9120 => "00111010", 9122 => "00101111", 9125 => "01001111", 9130 => "10010100", 9136 => "01010111", 9140 => "11010111", 9141 => "11000000", 9142 => "00011000", 9143 => "10001101", 9144 => "10110010", 9145 => "00001000", 9147 => "00000001", 9148 => "01111010", 9149 => "11110101", 9150 => "11011011", 9151 => "11010111", 9152 => "00010001", 9155 => "01001110", 9158 => "11100000", 9160 => "01110100", 9163 => "10101111", 9164 => "10011100", 9165 => "11011010", 9166 => "11101101", 9169 => "10011110", 9170 => "01110111", 9171 => "11101100", 9173 => "10100111", 9175 => "10011111", 9176 => "10100101", 9180 => "01011011", 9181 => "10101001", 9184 => "10011000", 9185 => "10100101", 9186 => "11110110", 9192 => "01001011", 9201 => "10001010", 9203 => "00011010", 9204 => "01001101", 9206 => "10000011", 9207 => "00010010", 9208 => "00011101", 9209 => "11010101", 9210 => "10010110", 9214 => "10100111", 9215 => "00100011", 9216 => "11110111", 9217 => "10000011", 9219 => "10111010", 9220 => "01001001", 9221 => "11111000", 9222 => "01111001", 9224 => "10011100", 9228 => "11101001", 9229 => "10010000", 9233 => "10100011", 9234 => "10000111", 9235 => "10011000", 9237 => "00110001", 9238 => "01001111", 9243 => "10011000", 9245 => "11111111", 9246 => "00000110", 9247 => "00010110", 9248 => "00101100", 9251 => "01000000", 9252 => "11001111", 9254 => "01101111", 9257 => "01101010", 9259 => "11010110", 9261 => "11100101", 9262 => "00110110", 9263 => "00111110", 9264 => "10001111", 9265 => "01100101", 9270 => "11010011", 9271 => "00101100", 9273 => "00101001", 9274 => "01000001", 9275 => "11110011", 9276 => "10001101", 9277 => "11111011", 9284 => "11011110", 9285 => "11010100", 9289 => "11001110", 9290 => "10001010", 9291 => "11010101", 9293 => "01000100", 9294 => "00100100", 9296 => "01110010", 9297 => "10011101", 9299 => "01100011", 9300 => "00100011", 9302 => "10101100", 9303 => "11110101", 9305 => "10111100", 9306 => "10111101", 9307 => "00010100", 9311 => "10001000", 9316 => "11110011", 9318 => "01110110", 9321 => "01010101", 9323 => "10011001", 9324 => "11101101", 9325 => "11110010", 9327 => "11001100", 9328 => "10010001", 9329 => "01000111", 9330 => "00100011", 9331 => "01101111", 9332 => "10101011", 9337 => "00101110", 9338 => "10110001", 9340 => "01000101", 9341 => "11000011", 9342 => "11010001", 9344 => "01100011", 9345 => "11010111", 9350 => "00000011", 9351 => "11110101", 9353 => "01100010", 9356 => "01101000", 9361 => "01110111", 9364 => "00100111", 9365 => "10001111", 9366 => "10011010", 9368 => "10010011", 9369 => "00011010", 9372 => "11111111", 9373 => "00000101", 9375 => "00110000", 9376 => "01100111", 9377 => "01111101", 9378 => "00111111", 9381 => "00110110", 9383 => "11111001", 9386 => "01010010", 9387 => "11001101", 9389 => "11011010", 9392 => "01011001", 9393 => "01011101", 9395 => "10101100", 9397 => "00111100", 9398 => "00101000", 9401 => "01111101", 9402 => "00101001", 9403 => "10100010", 9406 => "00101100", 9408 => "00011101", 9410 => "01011001", 9413 => "11000011", 9414 => "00111110", 9415 => "00110101", 9417 => "10010110", 9418 => "00000001", 9421 => "11010001", 9422 => "11001010", 9423 => "00100010", 9424 => "11101011", 9426 => "00011000", 9428 => "10111010", 9429 => "01011101", 9430 => "00001111", 9437 => "10100000", 9439 => "11011010", 9441 => "00000111", 9444 => "10000110", 9445 => "01010000", 9446 => "01001100", 9450 => "10001100", 9452 => "10111011", 9454 => "00010110", 9455 => "00110001", 9457 => "01011001", 9460 => "11110100", 9461 => "00011100", 9466 => "10011101", 9467 => "11001101", 9469 => "10110110", 9470 => "10110000", 9471 => "00111111", 9474 => "00011110", 9475 => "00010111", 9476 => "01001011", 9478 => "10011101", 9480 => "10100011", 9487 => "01010010", 9488 => "00011111", 9490 => "10100001", 9496 => "01101001", 9501 => "01010100", 9502 => "11101011", 9504 => "00101110", 9505 => "00110100", 9507 => "11010011", 9508 => "10000100", 9511 => "01111001", 9512 => "01100011", 9515 => "11010010", 9516 => "11011011", 9517 => "11101010", 9518 => "01000100", 9519 => "11100001", 9520 => "11011110", 9521 => "01100100", 9525 => "00000001", 9526 => "00010001", 9528 => "00011110", 9529 => "11110111", 9533 => "10100100", 9534 => "10011101", 9535 => "11011110", 9538 => "01111100", 9539 => "10111011", 9540 => "11001100", 9541 => "01111000", 9543 => "10101101", 9547 => "00101010", 9548 => "00010100", 9549 => "10110000", 9550 => "01001101", 9551 => "00110011", 9552 => "11011100", 9556 => "10111100", 9559 => "11000101", 9560 => "01011011", 9562 => "10100111", 9564 => "10101011", 9566 => "00000010", 9567 => "11111000", 9568 => "00110010", 9570 => "01111110", 9572 => "10000001", 9576 => "00100101", 9577 => "11110110", 9579 => "00111101", 9580 => "01001101", 9581 => "10101001", 9582 => "01000011", 9586 => "11100101", 9587 => "10100010", 9591 => "11100111", 9592 => "01001110", 9594 => "11101010", 9596 => "01101110", 9597 => "00100001", 9599 => "01000000", 9602 => "10101010", 9604 => "01100101", 9607 => "10100110", 9609 => "01000111", 9612 => "01110111", 9615 => "10001110", 9616 => "10000000", 9617 => "00010001", 9618 => "00111111", 9619 => "10110001", 9623 => "01011101", 9624 => "00111011", 9627 => "00100101", 9628 => "00001011", 9635 => "00010111", 9638 => "11010000", 9640 => "00010111", 9643 => "00000011", 9644 => "11000110", 9645 => "01110010", 9647 => "01000110", 9648 => "10011001", 9650 => "10001100", 9654 => "00101100", 9657 => "01100001", 9661 => "11000101", 9664 => "01111100", 9666 => "11111010", 9669 => "01001010", 9670 => "00100111", 9671 => "10101110", 9672 => "00010110", 9673 => "00111011", 9675 => "00101110", 9676 => "01100011", 9677 => "10010100", 9680 => "11111010", 9681 => "00111111", 9687 => "10010010", 9690 => "01100011", 9694 => "01101101", 9696 => "00100101", 9697 => "00110010", 9698 => "00011001", 9699 => "10100011", 9700 => "01011011", 9703 => "00010110", 9705 => "01110000", 9708 => "01000011", 9709 => "10011110", 9713 => "10010010", 9716 => "01001101", 9717 => "11101100", 9719 => "00101000", 9720 => "10000110", 9723 => "00001101", 9724 => "10000101", 9725 => "01101000", 9726 => "11011100", 9727 => "00000001", 9729 => "01111011", 9730 => "10010010", 9732 => "00101011", 9736 => "10001110", 9737 => "01001011", 9740 => "00100001", 9742 => "00010111", 9746 => "10011011", 9751 => "11110010", 9753 => "01100000", 9755 => "00010000", 9760 => "01110100", 9761 => "01000110", 9764 => "11000000", 9768 => "11010000", 9770 => "00001101", 9773 => "11101001", 9775 => "10111111", 9776 => "11100010", 9777 => "11001110", 9778 => "01110010", 9779 => "11111100", 9781 => "11011100", 9782 => "10011000", 9783 => "01001111", 9785 => "11000111", 9790 => "10010011", 9793 => "00100010", 9794 => "01100111", 9796 => "11101110", 9798 => "11101111", 9799 => "01100100", 9800 => "00010111", 9803 => "01000101", 9804 => "10111000", 9807 => "11011110", 9808 => "11101100", 9809 => "01010001", 9810 => "11110010", 9811 => "11110001", 9812 => "10100101", 9813 => "10111100", 9814 => "11100111", 9818 => "11011000", 9819 => "10111101", 9820 => "01010011", 9823 => "10100001", 9825 => "10111011", 9827 => "00101101", 9829 => "01101000", 9834 => "10011010", 9838 => "01111011", 9840 => "10111001", 9842 => "11101010", 9843 => "01010001", 9845 => "01110010", 9847 => "11000000", 9850 => "10001101", 9851 => "10001010", 9852 => "00011110", 9854 => "00001111", 9864 => "11000110", 9870 => "10000000", 9872 => "01000100", 9873 => "01100001", 9878 => "01110001", 9879 => "00011111", 9882 => "01001100", 9883 => "01101111", 9884 => "01101111", 9885 => "11010111", 9887 => "11111100", 9888 => "00111111", 9891 => "00001111", 9892 => "00110000", 9893 => "11111010", 9899 => "00010000", 9900 => "01001001", 9902 => "10111101", 9904 => "00010001", 9907 => "10011111", 9908 => "01111101", 9910 => "10100000", 9912 => "10010011", 9914 => "10001001", 9915 => "00000110", 9917 => "00110100", 9919 => "01010101", 9920 => "10100011", 9923 => "00101110", 9925 => "10110000", 9926 => "01100001", 9927 => "01111110", 9928 => "01010010", 9932 => "01110010", 9933 => "01100000", 9935 => "10010000", 9936 => "00111100", 9937 => "10110100", 9938 => "00100111", 9939 => "00100110", 9941 => "00101110", 9942 => "11011100", 9943 => "01111011", 9945 => "01001010", 9946 => "01001011", 9947 => "11011111", 9948 => "11110111", 9950 => "01000001", 9951 => "00000011", 9953 => "01001111", 9957 => "01011101", 9958 => "00001011", 9959 => "00001111", 9960 => "00111101", 9962 => "11010111", 9963 => "11001001", 9966 => "11101010", 9968 => "11010110", 9970 => "00000100", 9971 => "10010111", 9972 => "01100100", 9973 => "01010010", 9974 => "11100011", 9975 => "11011011", 9976 => "00001011", 9977 => "00111100", 9978 => "10110100", 9979 => "01101111", 9982 => "01000110", 9983 => "01100110", 9984 => "10111011", 9985 => "00010001", 9986 => "00100111", 9989 => "10110110", 9991 => "01000001", 9993 => "11111010", 9995 => "01011001", 9997 => "11001010", 9998 => "11111110", 10002 => "00111010", 10003 => "01110001", 10005 => "01111011", 10007 => "01001010", 10009 => "00001010", 10013 => "11111001", 10015 => "01100001", 10017 => "10101110", 10018 => "10110010", 10019 => "10100001", 10020 => "10011011", 10023 => "01110001", 10025 => "00001111", 10026 => "11100111", 10028 => "10011110", 10029 => "01011111", 10032 => "01101111", 10034 => "00110001", 10036 => "10100110", 10037 => "00011111", 10038 => "01011111", 10042 => "00100101", 10043 => "11111011", 10044 => "00111111", 10045 => "11111000", 10047 => "00110010", 10048 => "10000010", 10049 => "11110011", 10051 => "00101110", 10052 => "11000001", 10053 => "01111101", 10059 => "01001111", 10060 => "01011100", 10061 => "11110010", 10066 => "11000010", 10067 => "11010000", 10070 => "00011001", 10076 => "00001101", 10077 => "01111110", 10078 => "00001110", 10080 => "01001110", 10082 => "01110110", 10084 => "11100001", 10088 => "10111110", 10089 => "01101011", 10092 => "00001000", 10093 => "10110001", 10096 => "10110000", 10097 => "01101010", 10099 => "00111011", 10101 => "01110001", 10103 => "01100010", 10106 => "10110011", 10108 => "10011001", 10110 => "10101011", 10111 => "11000001", 10112 => "10010010", 10114 => "01100001", 10115 => "10010000", 10117 => "00001010", 10119 => "11000111", 10120 => "11000110", 10122 => "11001100", 10123 => "10100111", 10124 => "11101110", 10126 => "00110111", 10127 => "10111110", 10128 => "00011100", 10130 => "10011110", 10133 => "01001100", 10141 => "10000110", 10142 => "10111110", 10144 => "00111111", 10145 => "11111111", 10146 => "01010101", 10147 => "01000101", 10148 => "01001001", 10150 => "11010110", 10152 => "00100100", 10155 => "00011010", 10156 => "01101111", 10158 => "01010110", 10159 => "11011101", 10162 => "10111110", 10163 => "00000101", 10165 => "11110110", 10167 => "01010000", 10168 => "01111010", 10169 => "11011011", 10170 => "01000001", 10171 => "01000101", 10172 => "00111101", 10176 => "00110001", 10177 => "00100000", 10178 => "11011100", 10182 => "10100101", 10185 => "11110100", 10187 => "11011101", 10188 => "00010101", 10189 => "00011011", 10192 => "10111101", 10194 => "10111001", 10195 => "00101110", 10199 => "00100100", 10200 => "11010001", 10203 => "01101010", 10212 => "11010001", 10214 => "00110101", 10215 => "01000100", 10216 => "01111001", 10219 => "00011111", 10220 => "10010001", 10223 => "01100100", 10228 => "11110111", 10231 => "10010101", 10234 => "00111101", 10238 => "10100100", 10239 => "00100010", 10240 => "01111001", 10242 => "01011011", 10244 => "10101101", 10245 => "10000010", 10248 => "10010001", 10249 => "10101111", 10253 => "00001011", 10254 => "11001111", 10255 => "10111111", 10257 => "01110101", 10258 => "10110101", 10259 => "00100011", 10260 => "11000110", 10261 => "11111010", 10263 => "00110011", 10264 => "01100110", 10266 => "00011011", 10267 => "11010101", 10271 => "00000100", 10277 => "00001101", 10278 => "00001110", 10282 => "00010100", 10288 => "01110110", 10289 => "01100101", 10290 => "11010111", 10293 => "11100001", 10295 => "11001110", 10302 => "00011111", 10304 => "00101010", 10309 => "00110010", 10310 => "11011011", 10313 => "10111010", 10318 => "01100101", 10321 => "11010001", 10324 => "11110110", 10325 => "11000110", 10326 => "01001000", 10328 => "11101111", 10330 => "00100011", 10333 => "10011001", 10335 => "00101000", 10337 => "00000111", 10338 => "11111111", 10340 => "10001111", 10343 => "00000111", 10344 => "11010001", 10348 => "11001100", 10352 => "10101010", 10353 => "00011110", 10354 => "10100100", 10355 => "00100101", 10356 => "10101000", 10358 => "11011000", 10360 => "00000100", 10362 => "11101001", 10365 => "10001011", 10367 => "10010110", 10369 => "00010111", 10374 => "10101100", 10375 => "00100100", 10379 => "00001111", 10380 => "01100100", 10382 => "00111011", 10383 => "00000111", 10384 => "11100100", 10386 => "11100111", 10387 => "11110101", 10392 => "00110000", 10393 => "10100001", 10396 => "10011000", 10397 => "10011110", 10401 => "10000001", 10404 => "11011001", 10405 => "10011101", 10406 => "10100110", 10408 => "00011011", 10409 => "00001011", 10410 => "11100010", 10411 => "10000100", 10413 => "01011001", 10414 => "11011011", 10415 => "01111011", 10419 => "00011100", 10421 => "11010001", 10423 => "11100001", 10426 => "00100110", 10428 => "00111001", 10430 => "01101000", 10431 => "11010111", 10433 => "11001100", 10434 => "00010100", 10435 => "01111101", 10436 => "10011010", 10437 => "11010100", 10440 => "10100111", 10442 => "01110101", 10443 => "00011001", 10445 => "10110001", 10447 => "01111100", 10448 => "10010000", 10450 => "00111011", 10453 => "10101010", 10454 => "00100000", 10456 => "10101110", 10459 => "01010100", 10465 => "00110000", 10466 => "10010100", 10469 => "01000100", 10470 => "00010100", 10472 => "01101111", 10474 => "01110110", 10481 => "10000110", 10483 => "11111001", 10484 => "11010001", 10486 => "11100110", 10491 => "10110000", 10493 => "01010010", 10494 => "01000100", 10497 => "10101011", 10498 => "01100111", 10499 => "00001000", 10501 => "01011000", 10503 => "01111000", 10505 => "01000111", 10508 => "00010001", 10510 => "01101100", 10513 => "11000001", 10519 => "11000001", 10521 => "10110110", 10525 => "00101010", 10527 => "00011010", 10528 => "01001101", 10529 => "00100011", 10530 => "11001110", 10532 => "10011111", 10533 => "10001110", 10534 => "00000010", 10535 => "00011110", 10536 => "00010011", 10538 => "01111011", 10542 => "01110100", 10544 => "00010100", 10546 => "01000100", 10548 => "10001101", 10556 => "01100110", 10559 => "00101011", 10561 => "01110100", 10563 => "10000100", 10564 => "11100010", 10565 => "01010110", 10566 => "10001111", 10567 => "00100111", 10568 => "00011111", 10570 => "10101111", 10571 => "01010110", 10572 => "11110000", 10573 => "10101101", 10574 => "00000010", 10579 => "00100101", 10580 => "00011000", 10581 => "11110001", 10582 => "11110010", 10584 => "10110001", 10587 => "01010100", 10589 => "10010111", 10591 => "00110101", 10592 => "11000011", 10593 => "10001001", 10595 => "10101100", 10596 => "01001000", 10597 => "00001001", 10603 => "11001010", 10605 => "11111111", 10607 => "01101010", 10608 => "10010110", 10609 => "10101110", 10610 => "01110101", 10611 => "10000001", 10613 => "11111001", 10616 => "01101110", 10617 => "10100001", 10619 => "11111101", 10620 => "00101011", 10622 => "01000110", 10624 => "11100000", 10628 => "00001010", 10631 => "01011100", 10633 => "11001011", 10637 => "11000110", 10646 => "11100010", 10649 => "01111010", 10653 => "11001000", 10655 => "10011001", 10656 => "10110011", 10659 => "01011010", 10660 => "01111110", 10663 => "00110000", 10664 => "00101101", 10665 => "01100000", 10668 => "11000111", 10669 => "00010111", 10670 => "01111100", 10676 => "11100000", 10678 => "11000010", 10681 => "00111011", 10682 => "01010111", 10684 => "11110100", 10686 => "10101001", 10688 => "01000100", 10689 => "11001110", 10691 => "01011111", 10693 => "10100011", 10696 => "00011101", 10698 => "10110111", 10699 => "00010100", 10700 => "11010101", 10701 => "01110001", 10702 => "01111011", 10707 => "11011011", 10708 => "11110010", 10709 => "01100110", 10712 => "01010000", 10713 => "10111000", 10714 => "00100001", 10719 => "00111001", 10721 => "10101001", 10723 => "10100000", 10725 => "00010011", 10728 => "11110000", 10730 => "01011100", 10733 => "11011100", 10734 => "00010010", 10736 => "00011110", 10737 => "00010100", 10738 => "00001010", 10739 => "10110100", 10743 => "10100100", 10745 => "00101101", 10747 => "00100010", 10748 => "00100101", 10750 => "01111110", 10755 => "10010000", 10758 => "01100001", 10759 => "10100001", 10760 => "10001001", 10761 => "00000011", 10762 => "01110101", 10765 => "11000111", 10766 => "10011000", 10769 => "11111001", 10770 => "11010011", 10771 => "10100100", 10772 => "10000101", 10773 => "11010101", 10774 => "11110011", 10777 => "00010000", 10780 => "10101111", 10781 => "01101101", 10788 => "00100100", 10790 => "11001011", 10795 => "10001011", 10796 => "10010110", 10797 => "01011111", 10798 => "10001000", 10800 => "01001111", 10802 => "10001011", 10803 => "00011100", 10809 => "11001000", 10810 => "11001111", 10813 => "10110010", 10814 => "11010101", 10815 => "11000011", 10816 => "11110111", 10817 => "01101110", 10818 => "11110000", 10820 => "01000111", 10822 => "00001100", 10824 => "01000001", 10825 => "00101011", 10830 => "10001011", 10833 => "00010001", 10836 => "11000101", 10837 => "11111100", 10843 => "01111000", 10845 => "10011001", 10847 => "01101110", 10848 => "11011101", 10849 => "11001000", 10851 => "00111011", 10852 => "10010001", 10853 => "11010011", 10855 => "10110111", 10856 => "01001100", 10858 => "11111101", 10859 => "10001101", 10863 => "10000100", 10864 => "10110100", 10866 => "01010000", 10870 => "01010101", 10872 => "11011100", 10874 => "00001011", 10875 => "11101101", 10876 => "10011110", 10881 => "01001001", 10882 => "10100110", 10883 => "01100010", 10887 => "00011111", 10888 => "01111100", 10890 => "01000101", 10892 => "01011110", 10893 => "11001010", 10896 => "00101011", 10898 => "01010001", 10901 => "10011101", 10903 => "11110011", 10904 => "10010001", 10905 => "10101010", 10906 => "11100011", 10908 => "01001110", 10910 => "01001011", 10913 => "11111011", 10914 => "01001001", 10915 => "01110101", 10921 => "10100001", 10922 => "11100100", 10923 => "01101011", 10924 => "01100000", 10925 => "10001111", 10927 => "11100000", 10929 => "01011111", 10930 => "01100011", 10931 => "11000011", 10933 => "01111000", 10934 => "00101110", 10935 => "00101001", 10937 => "11111011", 10938 => "01011000", 10941 => "11011100", 10945 => "11110010", 10946 => "01100101", 10948 => "00010001", 10951 => "00010010", 10954 => "00101001", 10955 => "00111001", 10956 => "11110101", 10961 => "00110100", 10962 => "00101111", 10964 => "11000110", 10965 => "10110011", 10967 => "11000101", 10969 => "01001111", 10971 => "10001100", 10975 => "10000010", 10978 => "01010001", 10979 => "11111101", 10981 => "01100001", 10982 => "11011000", 10984 => "00001011", 10986 => "01010100", 10988 => "00101111", 10996 => "01101110", 10997 => "11111000", 10998 => "10101101", 11003 => "00001111", 11004 => "01000010", 11005 => "10010110", 11009 => "00100111", 11014 => "00101101", 11015 => "01011100", 11018 => "11100111", 11020 => "00011100", 11021 => "01100111", 11022 => "00111101", 11023 => "01000010", 11026 => "11101001", 11027 => "01111001", 11030 => "10100101", 11033 => "00011010", 11034 => "01011000", 11036 => "00100011", 11038 => "01101011", 11041 => "10101100", 11042 => "10111100", 11043 => "01110110", 11044 => "10001010", 11045 => "01010101", 11046 => "10110011", 11047 => "11011100", 11049 => "10010100", 11050 => "11000000", 11051 => "01101100", 11052 => "10001011", 11053 => "01100000", 11054 => "01011111", 11055 => "01110011", 11057 => "01010010", 11059 => "11110011", 11060 => "11100101", 11063 => "10111011", 11066 => "10100100", 11067 => "01000010", 11069 => "11010101", 11070 => "11101010", 11072 => "01101100", 11076 => "11011100", 11079 => "10000110", 11082 => "01111101", 11087 => "11001010", 11088 => "00011101", 11090 => "01101110", 11093 => "00101001", 11094 => "00000111", 11095 => "00011110", 11097 => "11110100", 11098 => "01111010", 11099 => "10110010", 11101 => "10110100", 11102 => "11101100", 11105 => "00100011", 11111 => "10111111", 11114 => "00010100", 11115 => "11011001", 11116 => "01100111", 11121 => "01010111", 11125 => "00101111", 11126 => "10001101", 11129 => "11010011", 11130 => "10011011", 11133 => "00011101", 11134 => "10000100", 11136 => "00000100", 11137 => "11110110", 11142 => "01011010", 11144 => "11110110", 11145 => "10001101", 11148 => "10110101", 11150 => "10100110", 11151 => "01100111", 11155 => "10101010", 11157 => "00101001", 11159 => "10000001", 11161 => "10100001", 11164 => "01001111", 11165 => "11111000", 11170 => "11101100", 11171 => "01111010", 11174 => "01011011", 11175 => "10011111", 11177 => "01000110", 11179 => "01011100", 11180 => "10100011", 11182 => "00100100", 11184 => "11111010", 11187 => "00010011", 11188 => "01100100", 11190 => "11011000", 11191 => "11111011", 11192 => "11000000", 11195 => "10010000", 11198 => "01111000", 11199 => "11011100", 11205 => "01000111", 11206 => "10100011", 11207 => "01101011", 11208 => "00101010", 11210 => "00111110", 11216 => "10010101", 11217 => "01010110", 11218 => "00000111", 11219 => "11010111", 11224 => "11110010", 11225 => "10100000", 11226 => "10100001", 11227 => "00100010", 11228 => "00111111", 11229 => "01111111", 11231 => "10001001", 11236 => "00110100", 11238 => "10000111", 11239 => "11001010", 11241 => "01110110", 11243 => "10010110", 11244 => "10101001", 11245 => "10101100", 11247 => "10111000", 11249 => "00101011", 11250 => "01110001", 11251 => "10000110", 11253 => "11010101", 11255 => "00010001", 11257 => "01001111", 11263 => "11001110", 11268 => "11011000", 11273 => "10100001", 11275 => "10111001", 11276 => "01110101", 11277 => "00100011", 11279 => "10011010", 11282 => "11001101", 11284 => "11101000", 11285 => "10011011", 11286 => "11010111", 11289 => "01000010", 11291 => "01010101", 11293 => "10010001", 11294 => "11001010", 11295 => "00011111", 11296 => "11011011", 11299 => "11100111", 11300 => "01111010", 11303 => "01000000", 11304 => "11010011", 11305 => "11011100", 11306 => "01110000", 11309 => "00101101", 11310 => "00010100", 11311 => "11101111", 11312 => "10000101", 11315 => "01111000", 11318 => "00000100", 11319 => "00011101", 11320 => "10100111", 11323 => "01011110", 11324 => "10110111", 11326 => "10011110", 11327 => "01001011", 11328 => "00101000", 11331 => "01110101", 11342 => "00110100", 11343 => "11011100", 11347 => "01101001", 11348 => "01101111", 11351 => "10010101", 11352 => "10011011", 11353 => "01101011", 11356 => "01011001", 11357 => "00011101", 11359 => "10111000", 11362 => "10100100", 11364 => "11010010", 11365 => "01001000", 11367 => "11001101", 11368 => "00110011", 11372 => "11011110", 11376 => "11010101", 11379 => "00011101", 11380 => "11110101", 11381 => "00100010", 11383 => "10010001", 11386 => "00101111", 11389 => "00011000", 11390 => "10010010", 11391 => "10100000", 11392 => "10110000", 11395 => "01110111", 11396 => "00111010", 11397 => "00111000", 11398 => "11100100", 11399 => "00111100", 11402 => "00001100", 11403 => "01110000", 11404 => "01110101", 11405 => "11011011", 11406 => "01111101", 11407 => "10001110", 11409 => "11001001", 11411 => "11110101", 11413 => "11110101", 11414 => "00011001", 11415 => "11000111", 11416 => "10111001", 11417 => "11100110", 11418 => "01110000", 11419 => "11100110", 11420 => "01001111", 11421 => "00001100", 11422 => "10100000", 11425 => "10100111", 11427 => "10110101", 11429 => "11100100", 11431 => "00100101", 11433 => "11011101", 11436 => "01110110", 11437 => "10100000", 11439 => "10101011", 11440 => "10101010", 11441 => "01001100", 11442 => "01110100", 11443 => "01111001", 11444 => "11101110", 11446 => "00010001", 11448 => "10110100", 11449 => "00111101", 11451 => "11000011", 11452 => "10101000", 11453 => "10001011", 11454 => "00110011", 11456 => "00011001", 11460 => "10100110", 11462 => "11111110", 11464 => "10011100", 11466 => "01000000", 11467 => "11101001", 11470 => "00100100", 11473 => "01110110", 11477 => "01011110", 11478 => "11001001", 11479 => "10111000", 11481 => "10101010", 11482 => "11100000", 11483 => "00101100", 11485 => "10100010", 11488 => "10000010", 11489 => "00100000", 11491 => "11111011", 11493 => "01011001", 11497 => "00110001", 11499 => "00110000", 11502 => "11001001", 11505 => "00010110", 11509 => "00111000", 11513 => "11111010", 11517 => "01111001", 11520 => "10000111", 11524 => "10111000", 11529 => "11111011", 11535 => "10101001", 11538 => "11111010", 11539 => "10011010", 11540 => "01101110", 11543 => "01010011", 11546 => "11000001", 11550 => "01001000", 11551 => "10111000", 11554 => "11101110", 11558 => "10000010", 11559 => "10101101", 11560 => "10111000", 11561 => "01011011", 11562 => "11111010", 11565 => "11101100", 11569 => "10100111", 11573 => "01001011", 11574 => "10001101", 11580 => "01010110", 11581 => "01110111", 11582 => "01111111", 11586 => "00010001", 11589 => "00110100", 11592 => "00010111", 11596 => "11001010", 11597 => "10100100", 11599 => "00101011", 11601 => "00101101", 11602 => "01110001", 11604 => "00101011", 11605 => "11011101", 11608 => "01001010", 11609 => "11110000", 11611 => "00111101", 11613 => "00101101", 11614 => "00010001", 11615 => "00110110", 11618 => "10011100", 11620 => "01010101", 11621 => "10001011", 11623 => "00000010", 11625 => "11101111", 11628 => "11110000", 11629 => "00110111", 11630 => "01111111", 11636 => "01011010", 11640 => "10101101", 11642 => "00100100", 11645 => "11100101", 11649 => "11110110", 11651 => "01010011", 11656 => "00010000", 11660 => "00110111", 11661 => "00011110", 11663 => "00011001", 11664 => "11010001", 11667 => "10101110", 11668 => "01100001", 11669 => "01010100", 11672 => "10100001", 11676 => "11001111", 11678 => "01000100", 11680 => "00101000", 11684 => "01010100", 11687 => "00010111", 11688 => "10110000", 11690 => "11110001", 11691 => "01011000", 11692 => "01010010", 11693 => "00111101", 11694 => "10110010", 11695 => "01011000", 11696 => "10111001", 11697 => "10110100", 11700 => "01101001", 11704 => "11100100", 11705 => "01001100", 11706 => "00101101", 11707 => "10011001", 11709 => "01111001", 11710 => "01110000", 11711 => "11010010", 11713 => "00000001", 11714 => "01011100", 11715 => "00001101", 11720 => "00101001", 11721 => "01110111", 11723 => "00000101", 11724 => "01100000", 11731 => "01001000", 11732 => "10001111", 11733 => "10010100", 11734 => "00111010", 11736 => "01101010", 11739 => "11101111", 11741 => "11101111", 11743 => "10111011", 11744 => "01100010", 11748 => "11111100", 11750 => "01010001", 11751 => "10011010", 11754 => "10000101", 11755 => "11000000", 11759 => "10001011", 11761 => "00011000", 11762 => "10110101", 11764 => "00110111", 11765 => "01101010", 11766 => "10000001", 11767 => "11011010", 11768 => "10100001", 11771 => "10100000", 11776 => "01001011", 11777 => "10010110", 11778 => "10100111", 11779 => "10000010", 11782 => "01001000", 11785 => "11000111", 11791 => "11110111", 11794 => "11001011", 11795 => "10011101", 11796 => "11011001", 11802 => "01010001", 11807 => "01011001", 11809 => "11001011", 11810 => "10110111", 11811 => "10101111", 11814 => "11100000", 11816 => "01000100", 11819 => "01110100", 11821 => "11001011", 11828 => "11010110", 11829 => "00000011", 11831 => "01010100", 11832 => "00001100", 11839 => "01110000", 11840 => "00100110", 11841 => "00110000", 11843 => "11000010", 11851 => "10010110", 11853 => "00111101", 11855 => "01010000", 11857 => "01000010", 11859 => "00001100", 11860 => "00101000", 11861 => "11011110", 11862 => "00100101", 11863 => "11011010", 11865 => "10101011", 11868 => "11110001", 11869 => "11111001", 11870 => "01001100", 11871 => "11011111", 11874 => "01011111", 11877 => "10111010", 11878 => "11110001", 11879 => "10111110", 11880 => "10101000", 11881 => "10011010", 11885 => "01111101", 11887 => "10111110", 11888 => "11000110", 11891 => "00111101", 11895 => "01100110", 11901 => "11010011", 11908 => "11101001", 11911 => "10101010", 11912 => "01011100", 11915 => "11000101", 11916 => "10000100", 11917 => "00111111", 11918 => "10000110", 11924 => "10101001", 11926 => "10000100", 11927 => "01000001", 11928 => "11100100", 11931 => "11001101", 11933 => "10010010", 11935 => "11101111", 11937 => "11011101", 11938 => "01110000", 11939 => "10100111", 11940 => "00001000", 11944 => "01110000", 11945 => "00000001", 11946 => "11000110", 11952 => "01111011", 11954 => "00101111", 11956 => "11101100", 11959 => "01111010", 11960 => "01010011", 11961 => "10100111", 11962 => "10000000", 11963 => "01001010", 11965 => "10011111", 11967 => "11100110", 11972 => "00011011", 11975 => "01111000", 11978 => "00010001", 11982 => "00000111", 11984 => "10001000", 11987 => "01011011", 11992 => "01111110", 11994 => "00000110", 11995 => "11000000", 12000 => "00101110", 12003 => "00111011", 12004 => "00110101", 12005 => "10111110", 12006 => "01011000", 12007 => "11101001", 12010 => "00010100", 12011 => "10101011", 12012 => "01111000", 12013 => "11001000", 12015 => "11110111", 12017 => "00001101", 12018 => "10010010", 12019 => "00011011", 12020 => "00100000", 12022 => "10011111", 12027 => "01011110", 12028 => "10000011", 12033 => "11111010", 12040 => "10010011", 12042 => "10000111", 12043 => "00101110", 12045 => "00110011", 12048 => "11100001", 12050 => "11101010", 12053 => "11101100", 12055 => "01100100", 12057 => "10110001", 12060 => "01101011", 12062 => "11110111", 12064 => "10000111", 12067 => "00111001", 12068 => "11011111", 12071 => "10000111", 12072 => "01011000", 12076 => "11000000", 12078 => "01001000", 12082 => "01101010", 12084 => "10010001", 12088 => "10000011", 12089 => "11111101", 12090 => "00100001", 12093 => "00101111", 12095 => "01110110", 12096 => "00101101", 12104 => "11010101", 12105 => "00000110", 12106 => "11111111", 12107 => "11101010", 12109 => "11011001", 12111 => "00110100", 12113 => "01111101", 12114 => "01101000", 12116 => "01010011", 12119 => "01011011", 12120 => "10000100", 12121 => "01000010", 12123 => "11010111", 12124 => "11011011", 12126 => "00111000", 12129 => "10000110", 12132 => "00011011", 12136 => "10001011", 12138 => "01001011", 12140 => "10110011", 12141 => "11100111", 12142 => "01010101", 12143 => "11001011", 12149 => "00111001", 12153 => "10011011", 12161 => "10001011", 12165 => "01010010", 12167 => "00000111", 12170 => "11000011", 12172 => "01010100", 12174 => "10101101", 12175 => "10100100", 12179 => "11100001", 12188 => "11011010", 12189 => "01001011", 12190 => "11000110", 12191 => "01101011", 12198 => "11000001", 12202 => "11101000", 12209 => "10100111", 12211 => "00010110", 12213 => "01000000", 12214 => "11001100", 12215 => "10111010", 12216 => "11100111", 12217 => "10001001", 12220 => "01000001", 12222 => "00111001", 12223 => "11010100", 12224 => "00101101", 12227 => "00111001", 12228 => "00101100", 12229 => "11010010", 12232 => "11000001", 12235 => "01101000", 12236 => "01000010", 12238 => "10010110", 12240 => "01110000", 12241 => "11111000", 12242 => "01001011", 12243 => "01000101", 12246 => "10110110", 12247 => "00000111", 12248 => "10011100", 12249 => "10010011", 12250 => "10110100", 12254 => "01100010", 12260 => "01001100", 12261 => "01100011", 12262 => "01011101", 12263 => "10111011", 12265 => "01010110", 12267 => "10000101", 12268 => "01100000", 12269 => "10000011", 12271 => "11000111", 12272 => "00001110", 12275 => "01100001", 12280 => "01100010", 12281 => "01100000", 12285 => "11101001", 12288 => "10110110", 12289 => "00001110", 12291 => "11100000", 12293 => "11111000", 12294 => "00001010", 12297 => "10110101", 12300 => "10000010", 12302 => "10110011", 12303 => "11011001", 12306 => "01010001", 12307 => "00111010", 12309 => "11001101", 12310 => "10111110", 12311 => "01100011", 12313 => "01001001", 12314 => "11101110", 12317 => "00011001", 12318 => "11111000", 12319 => "10110101", 12320 => "10100010", 12321 => "11010010", 12322 => "10010010", 12324 => "00011001", 12325 => "01001110", 12326 => "00001011", 12328 => "00011111", 12329 => "11101001", 12330 => "11110011", 12331 => "01010100", 12332 => "00111010", 12333 => "01111110", 12334 => "00010010", 12335 => "01010001", 12336 => "00101100", 12340 => "00011111", 12341 => "10010000", 12344 => "10111001", 12348 => "00101101", 12353 => "00011010", 12354 => "00110001", 12355 => "01010011", 12356 => "11101101", 12357 => "10011111", 12360 => "01101001", 12362 => "11001111", 12365 => "11011010", 12369 => "11001100", 12370 => "01011000", 12372 => "00100001", 12374 => "01100111", 12375 => "11000011", 12376 => "01100000", 12379 => "11100101", 12381 => "11010000", 12384 => "00110010", 12388 => "01111111", 12395 => "11100100", 12396 => "11010010", 12399 => "11000011", 12400 => "11110111", 12401 => "01001010", 12402 => "11011001", 12403 => "10100011", 12405 => "01010010", 12406 => "11100101", 12410 => "00100110", 12415 => "01100001", 12418 => "11010010", 12420 => "11000110", 12421 => "10110010", 12422 => "01110111", 12423 => "11011001", 12424 => "10010010", 12426 => "01101000", 12427 => "00011111", 12428 => "10010010", 12429 => "00100100", 12432 => "00001110", 12433 => "00001001", 12435 => "11110111", 12436 => "11100010", 12437 => "11101011", 12441 => "11110001", 12442 => "11110001", 12445 => "00101001", 12446 => "00100101", 12449 => "01110000", 12454 => "00010010", 12455 => "00010010", 12457 => "00101001", 12459 => "10110011", 12461 => "00111110", 12464 => "10011010", 12466 => "01111100", 12467 => "00001110", 12468 => "10111011", 12471 => "00101000", 12473 => "10001011", 12475 => "11110001", 12476 => "11101100", 12477 => "00110001", 12478 => "10011011", 12481 => "01100011", 12485 => "01100010", 12487 => "10011111", 12488 => "01011010", 12492 => "00001001", 12493 => "01101110", 12494 => "00100000", 12496 => "01110100", 12498 => "10000110", 12499 => "01100111", 12501 => "11011101", 12505 => "10100100", 12507 => "11011000", 12509 => "11110000", 12510 => "00000001", 12514 => "00110111", 12515 => "01110010", 12516 => "11100000", 12517 => "01111011", 12520 => "01011010", 12523 => "11011101", 12524 => "01110000", 12525 => "11110000", 12526 => "11000000", 12528 => "11011101", 12529 => "01000101", 12533 => "11011111", 12534 => "00110101", 12537 => "00100011", 12538 => "01110111", 12539 => "01000011", 12540 => "01101011", 12542 => "00101011", 12543 => "00000100", 12544 => "10000010", 12550 => "00100111", 12551 => "01011110", 12552 => "01111111", 12554 => "10000011", 12555 => "01100110", 12556 => "01011010", 12557 => "11011000", 12559 => "00001001", 12560 => "10110011", 12562 => "00011110", 12564 => "01101110", 12567 => "00011001", 12568 => "11100001", 12571 => "01111000", 12573 => "11011111", 12576 => "00011111", 12577 => "00001100", 12578 => "01110100", 12579 => "00011110", 12581 => "10111010", 12582 => "10000100", 12583 => "10100001", 12584 => "00110110", 12589 => "10100101", 12590 => "11111010", 12591 => "10001111", 12592 => "00100111", 12593 => "01110010", 12594 => "00001001", 12595 => "00111001", 12596 => "11111110", 12599 => "11010100", 12600 => "00010100", 12603 => "01001011", 12604 => "01111110", 12605 => "01000111", 12607 => "00101110", 12611 => "00010010", 12613 => "10110101", 12615 => "11010001", 12617 => "01100101", 12618 => "11110001", 12620 => "11000101", 12622 => "00111110", 12623 => "10111000", 12624 => "01111111", 12626 => "11000100", 12627 => "10001011", 12630 => "00110100", 12632 => "01001000", 12636 => "00110010", 12641 => "10010011", 12646 => "10100101", 12650 => "00001000", 12653 => "10101010", 12655 => "00001111", 12656 => "01100101", 12657 => "10100101", 12659 => "11111110", 12660 => "00100010", 12668 => "11010110", 12669 => "01100001", 12670 => "01011101", 12671 => "10111100", 12673 => "00110011", 12674 => "11000010", 12675 => "00101011", 12676 => "01111010", 12678 => "00110100", 12679 => "11001000", 12681 => "01011011", 12682 => "01101101", 12683 => "00101111", 12684 => "11101111", 12691 => "00100011", 12693 => "11001001", 12694 => "11011000", 12700 => "10011101", 12703 => "01000110", 12704 => "01010111", 12706 => "10110000", 12708 => "01011101", 12710 => "10100100", 12712 => "11101100", 12713 => "01100011", 12717 => "11000000", 12719 => "01110101", 12720 => "00100111", 12721 => "01101001", 12724 => "00001000", 12725 => "01011001", 12728 => "11100111", 12729 => "01011110", 12734 => "10001001", 12735 => "00011011", 12736 => "10000011", 12739 => "01000001", 12741 => "10100011", 12742 => "01110011", 12744 => "11000111", 12745 => "10011001", 12746 => "00011111", 12749 => "10100100", 12750 => "00010110", 12751 => "11101000", 12754 => "11010000", 12757 => "11110001", 12759 => "10101000", 12763 => "00101110", 12764 => "10110110", 12768 => "00111111", 12771 => "00000101", 12775 => "01110100", 12776 => "00110111", 12780 => "11010000", 12781 => "10000011", 12782 => "11100100", 12783 => "10010110", 12796 => "01111111", 12803 => "10000101", 12806 => "11001010", 12808 => "01101111", 12811 => "11000001", 12813 => "00010100", 12814 => "00110111", 12815 => "00001101", 12816 => "01001010", 12817 => "01001001", 12818 => "11110010", 12820 => "01010000", 12822 => "01011001", 12826 => "00010011", 12827 => "10001110", 12832 => "01011101", 12833 => "11001101", 12834 => "00000101", 12836 => "10110010", 12838 => "10100011", 12839 => "01111110", 12842 => "10011000", 12844 => "11011000", 12845 => "01100111", 12846 => "10100100", 12849 => "11001010", 12851 => "01011010", 12852 => "01110011", 12855 => "01111111", 12856 => "11101100", 12858 => "00000100", 12861 => "10001101", 12862 => "11011011", 12864 => "01000011", 12867 => "00011001", 12870 => "11010011", 12871 => "01011000", 12874 => "01100000", 12875 => "01010100", 12876 => "10110010", 12885 => "10001111", 12886 => "11100110", 12890 => "01100001", 12891 => "10110011", 12893 => "00100011", 12897 => "00010010", 12905 => "00000001", 12907 => "10110011", 12908 => "11101111", 12910 => "11010000", 12911 => "01111101", 12912 => "00000001", 12913 => "00000101", 12918 => "01110000", 12919 => "00001101", 12920 => "01110010", 12922 => "01011111", 12924 => "01011001", 12925 => "01011011", 12926 => "00101011", 12928 => "10101010", 12929 => "10100011", 12930 => "00100011", 12932 => "01000001", 12934 => "01010111", 12935 => "01010000", 12938 => "00101000", 12939 => "11000111", 12941 => "10001000", 12944 => "11111011", 12946 => "00000110", 12947 => "10111011", 12949 => "01001111", 12953 => "00010011", 12956 => "11101110", 12957 => "11110011", 12959 => "00101010", 12960 => "00101100", 12961 => "11000101", 12967 => "01111001", 12968 => "10101110", 12969 => "00100101", 12970 => "10001000", 12972 => "10010101", 12974 => "00001101", 12976 => "10001100", 12977 => "11110000", 12979 => "10110011", 12980 => "01111000", 12982 => "01011000", 12983 => "10010011", 12986 => "00010010", 12988 => "11101011", 12991 => "01011101", 12992 => "00010001", 12994 => "01000001", 12997 => "10001001", 13000 => "10001100", 13005 => "00100001", 13007 => "11010011", 13008 => "01000110", 13009 => "10101101", 13012 => "00101100", 13013 => "01011100", 13016 => "10010100", 13018 => "01110101", 13020 => "11110010", 13021 => "11001011", 13022 => "00101111", 13027 => "01100110", 13031 => "11111111", 13034 => "11010111", 13035 => "00111101", 13037 => "10101111", 13039 => "10001001", 13040 => "11001000", 13042 => "11101000", 13044 => "00110000", 13046 => "11100100", 13050 => "00001111", 13052 => "10000011", 13054 => "01011001", 13055 => "00010000", 13056 => "01110000", 13061 => "01010000", 13063 => "11110011", 13065 => "10010111", 13068 => "10110101", 13070 => "00011010", 13073 => "11001101", 13075 => "10010011", 13078 => "10010000", 13079 => "01010000", 13081 => "01100011", 13082 => "10011010", 13084 => "11001011", 13085 => "01100100", 13086 => "11000011", 13089 => "00110100", 13091 => "11101101", 13093 => "00110101", 13094 => "10001101", 13095 => "00101010", 13098 => "01000101", 13099 => "01111101", 13100 => "00000001", 13101 => "10010100", 13104 => "11011110", 13108 => "01110000", 13109 => "10101010", 13110 => "10001100", 13111 => "10100100", 13114 => "01000001", 13115 => "11000111", 13121 => "10100010", 13122 => "11111110", 13123 => "10100011", 13124 => "10011100", 13125 => "00011001", 13126 => "11001110", 13128 => "00111111", 13131 => "11000100", 13133 => "10110110", 13134 => "00101010", 13136 => "11001001", 13137 => "00110011", 13140 => "00010110", 13141 => "00100100", 13142 => "01001101", 13143 => "11100100", 13147 => "00001000", 13148 => "01001000", 13149 => "00111010", 13157 => "11111111", 13159 => "01000000", 13164 => "01111101", 13165 => "01010100", 13166 => "01011011", 13167 => "11000010", 13170 => "00100001", 13171 => "10001111", 13173 => "11001011", 13179 => "00110110", 13183 => "00100101", 13185 => "00001110", 13187 => "10010000", 13190 => "10110111", 13191 => "01110000", 13192 => "10100011", 13195 => "01100011", 13196 => "00011000", 13197 => "11001101", 13198 => "00111101", 13200 => "10101111", 13202 => "01010100", 13206 => "01110011", 13207 => "10011100", 13208 => "00001010", 13209 => "01100010", 13214 => "01000101", 13216 => "10100100", 13217 => "11010011", 13219 => "11010001", 13221 => "10110110", 13222 => "00000011", 13224 => "01000010", 13227 => "00010000", 13229 => "10000000", 13230 => "10110010", 13231 => "00101110", 13233 => "10011100", 13234 => "11000011", 13235 => "00001001", 13238 => "01111101", 13241 => "11001111", 13242 => "01011010", 13244 => "01001110", 13248 => "00010100", 13249 => "01001000", 13252 => "00010110", 13255 => "11011110", 13256 => "11011001", 13257 => "11000110", 13259 => "00110101", 13260 => "10011000", 13261 => "11111101", 13262 => "00111111", 13263 => "00101111", 13265 => "00011101", 13266 => "01000001", 13267 => "01101100", 13268 => "01001101", 13269 => "01011000", 13271 => "11000111", 13272 => "00111100", 13273 => "10110001", 13275 => "00000101", 13276 => "00110111", 13277 => "10110010", 13278 => "10100000", 13279 => "10101111", 13280 => "11101011", 13281 => "00101111", 13284 => "11101000", 13285 => "00010011", 13286 => "10101010", 13287 => "10101010", 13290 => "00000111", 13291 => "01101011", 13292 => "00101010", 13293 => "01000010", 13294 => "00101101", 13298 => "11111001", 13299 => "11010111", 13300 => "10000001", 13301 => "00111101", 13302 => "00110111", 13304 => "01001100", 13307 => "01101110", 13309 => "10000001", 13311 => "01100101", 13313 => "01100010", 13314 => "01111101", 13315 => "10011000", 13316 => "01001111", 13318 => "10111100", 13319 => "11110001", 13320 => "11101101", 13322 => "00111010", 13323 => "01010101", 13324 => "10001010", 13326 => "00011100", 13327 => "00110000", 13328 => "10110010", 13330 => "10011000", 13333 => "00101010", 13334 => "10011001", 13335 => "00001111", 13341 => "01110011", 13342 => "00100110", 13345 => "10010010", 13347 => "00010001", 13348 => "01000101", 13349 => "10001100", 13350 => "10001111", 13352 => "10111011", 13354 => "00010111", 13357 => "11100000", 13358 => "00100011", 13361 => "11100001", 13366 => "01110101", 13371 => "01100111", 13373 => "00111100", 13374 => "00011100", 13376 => "00111110", 13378 => "01111011", 13380 => "00001100", 13383 => "01110000", 13384 => "01101100", 13386 => "11010011", 13387 => "00001101", 13388 => "11110111", 13389 => "10001111", 13392 => "11000100", 13393 => "01101101", 13395 => "01100001", 13397 => "01010111", 13403 => "00100001", 13408 => "11101111", 13410 => "00100111", 13411 => "01000111", 13412 => "01000110", 13413 => "10001101", 13414 => "11001111", 13419 => "11110100", 13420 => "01111001", 13421 => "00111101", 13422 => "01111010", 13424 => "10001101", 13427 => "11011101", 13430 => "01001001", 13431 => "11010010", 13432 => "01010010", 13433 => "00010101", 13434 => "01010011", 13435 => "11011100", 13436 => "11110101", 13437 => "01100000", 13439 => "00010110", 13440 => "01000100", 13443 => "10100111", 13446 => "01100010", 13447 => "01101111", 13448 => "01011000", 13449 => "01101100", 13452 => "00001000", 13453 => "11111001", 13455 => "10010001", 13456 => "01100100", 13459 => "10011000", 13462 => "00011111", 13464 => "01111101", 13466 => "00000011", 13467 => "11010000", 13469 => "01110000", 13470 => "11101101", 13471 => "11001100", 13474 => "01100010", 13476 => "00111110", 13478 => "00001101", 13479 => "00110100", 13482 => "10110110", 13483 => "01110000", 13487 => "11111110", 13488 => "01101011", 13497 => "11001010", 13498 => "10010111", 13499 => "00000110", 13500 => "11001111", 13501 => "11001011", 13503 => "10110110", 13507 => "01101011", 13510 => "01110000", 13511 => "11000110", 13512 => "11100100", 13513 => "01010101", 13515 => "11110010", 13518 => "01000110", 13519 => "00110110", 13521 => "01101110", 13522 => "10110010", 13524 => "01011010", 13526 => "00110100", 13527 => "00101000", 13533 => "01111110", 13536 => "00001000", 13537 => "11000010", 13538 => "10000011", 13540 => "00101101", 13542 => "10011111", 13545 => "11000111", 13547 => "00111101", 13548 => "00100110", 13552 => "00011000", 13553 => "01101100", 13554 => "11101011", 13557 => "01010001", 13558 => "01000001", 13560 => "10011011", 13561 => "11000011", 13562 => "01000110", 13563 => "11101100", 13564 => "01111110", 13565 => "01100101", 13566 => "10100001", 13567 => "10111010", 13568 => "10111001", 13572 => "11101110", 13573 => "01011001", 13575 => "11100011", 13576 => "00110000", 13577 => "10010000", 13579 => "00100111", 13580 => "01000101", 13581 => "11101110", 13584 => "11010010", 13585 => "01101111", 13586 => "00111000", 13587 => "11000001", 13588 => "10101010", 13589 => "01111100", 13590 => "00010110", 13592 => "10010100", 13593 => "11001010", 13596 => "01000001", 13597 => "00011111", 13603 => "01101010", 13604 => "01010001", 13607 => "00010001", 13609 => "10110100", 13611 => "11001101", 13612 => "10000000", 13613 => "11001000", 13616 => "00011101", 13617 => "00101001", 13619 => "10010101", 13621 => "01111011", 13626 => "00100110", 13627 => "10000001", 13628 => "10101100", 13629 => "01101110", 13631 => "10111111", 13632 => "10010101", 13636 => "11001101", 13642 => "01111100", 13643 => "01000100", 13644 => "00100001", 13645 => "01010001", 13646 => "00010000", 13647 => "10011111", 13648 => "10111100", 13649 => "01011011", 13652 => "01011111", 13655 => "01010001", 13657 => "00100001", 13658 => "00111111", 13660 => "11111110", 13661 => "01010100", 13662 => "11010011", 13664 => "10110110", 13665 => "00010011", 13666 => "10000101", 13667 => "00110101", 13670 => "11101010", 13671 => "01110001", 13673 => "10101000", 13677 => "00001011", 13678 => "01011110", 13679 => "01100101", 13680 => "01000011", 13681 => "11110011", 13683 => "01111001", 13687 => "11000100", 13690 => "01010101", 13692 => "11010011", 13694 => "10110110", 13699 => "11101101", 13700 => "10110100", 13701 => "00010010", 13704 => "10000101", 13705 => "11111011", 13707 => "01001101", 13709 => "11111110", 13710 => "00100110", 13712 => "00011110", 13719 => "11110100", 13720 => "11111011", 13721 => "10000010", 13722 => "10110101", 13723 => "01100111", 13725 => "01110010", 13728 => "01000001", 13731 => "10101010", 13732 => "10011101", 13734 => "00110011", 13736 => "11010000", 13737 => "00110000", 13745 => "00010001", 13746 => "11000011", 13747 => "01011110", 13748 => "10010111", 13750 => "00010010", 13754 => "00111000", 13756 => "11110100", 13757 => "00110000", 13760 => "10101000", 13762 => "00001111", 13763 => "10010100", 13766 => "10110100", 13767 => "01101001", 13769 => "11011010", 13770 => "00010111", 13772 => "10111110", 13773 => "00111000", 13774 => "01000111", 13775 => "00110100", 13777 => "01001011", 13779 => "11100010", 13787 => "01011101", 13788 => "11010100", 13790 => "11000111", 13794 => "11101011", 13795 => "10110101", 13798 => "10000110", 13800 => "01110010", 13801 => "00010000", 13802 => "10011001", 13803 => "11100110", 13805 => "10110001", 13809 => "00001011", 13810 => "11011111", 13811 => "01101101", 13815 => "10111111", 13817 => "00110100", 13822 => "00100010", 13825 => "11000111", 13826 => "11111001", 13828 => "01100111", 13832 => "11010100", 13834 => "10111100", 13835 => "00111110", 13836 => "01000110", 13837 => "01110110", 13840 => "11001000", 13845 => "01101000", 13852 => "11001101", 13853 => "00111111", 13855 => "10010000", 13856 => "10010011", 13859 => "10001011", 13860 => "01111010", 13864 => "00111111", 13865 => "00000100", 13866 => "01111110", 13868 => "11111111", 13869 => "00011011", 13871 => "10101110", 13874 => "01101100", 13876 => "01111000", 13877 => "01010101", 13882 => "01110100", 13883 => "11010011", 13884 => "00011000", 13888 => "11101011", 13891 => "10010100", 13893 => "11111100", 13896 => "10001111", 13901 => "00110111", 13905 => "01100111", 13906 => "00010111", 13907 => "00111001", 13914 => "01111101", 13917 => "00100100", 13919 => "10001010", 13922 => "10111111", 13923 => "11011011", 13924 => "11000100", 13926 => "10000110", 13928 => "10100001", 13929 => "11001101", 13930 => "01011000", 13932 => "11001100", 13933 => "01111010", 13934 => "01101100", 13935 => "01111110", 13936 => "11010011", 13940 => "01000001", 13941 => "11100100", 13946 => "11000100", 13951 => "10011101", 13953 => "01110101", 13956 => "01010101", 13958 => "01111010", 13959 => "00001110", 13960 => "10011001", 13961 => "10101001", 13963 => "01010010", 13965 => "10001010", 13967 => "00100001", 13968 => "01110101", 13970 => "11110011", 13973 => "10010001", 13976 => "11100011", 13978 => "11011100", 13979 => "00000011", 13980 => "10010100", 13982 => "11001111", 13983 => "00001011", 13984 => "01001100", 13987 => "10000110", 13991 => "11111001", 13994 => "00011111", 13995 => "01010101", 13997 => "01101110", 13998 => "00111100", 14000 => "10011101", 14007 => "01111011", 14008 => "00011010", 14009 => "11011001", 14010 => "11101011", 14012 => "01011111", 14013 => "11011111", 14014 => "10100100", 14016 => "00100001", 14017 => "01110100", 14020 => "00000100", 14023 => "11110000", 14025 => "01000001", 14027 => "10110000", 14028 => "11100101", 14030 => "11001011", 14031 => "00011011", 14033 => "01010000", 14035 => "01111101", 14037 => "11101011", 14039 => "11100100", 14040 => "01001100", 14042 => "01010100", 14046 => "00001001", 14048 => "01111110", 14050 => "00001100", 14051 => "01110101", 14052 => "00010111", 14053 => "01010011", 14054 => "11100001", 14055 => "01111100", 14056 => "10110101", 14057 => "00111100", 14058 => "11010100", 14061 => "00000011", 14065 => "00100011", 14066 => "01010000", 14067 => "10011101", 14070 => "11010100", 14071 => "11010010", 14072 => "00111001", 14073 => "01001000", 14076 => "00010111", 14077 => "00110100", 14078 => "01100011", 14079 => "01010111", 14082 => "10001000", 14085 => "11101110", 14086 => "01100000", 14087 => "10001011", 14088 => "10000100", 14090 => "01110111", 14091 => "01100110", 14092 => "01110000", 14094 => "10001010", 14099 => "00110111", 14102 => "01101101", 14103 => "11001110", 14104 => "10001010", 14105 => "11101001", 14106 => "00100001", 14108 => "00101011", 14117 => "00110110", 14118 => "01110110", 14119 => "00011001", 14120 => "01111111", 14124 => "10010110", 14125 => "11110011", 14126 => "00100101", 14129 => "10111101", 14130 => "11101111", 14131 => "11110101", 14134 => "00010100", 14135 => "01111110", 14144 => "00111100", 14145 => "01011100", 14146 => "11011111", 14151 => "00010001", 14154 => "01100100", 14155 => "11111001", 14156 => "11010010", 14157 => "11101011", 14161 => "10100101", 14162 => "00101111", 14163 => "00101110", 14164 => "11010001", 14165 => "00100101", 14166 => "11010000", 14172 => "01111010", 14174 => "11011011", 14175 => "10000001", 14177 => "00101010", 14179 => "01010110", 14180 => "00100011", 14182 => "00110111", 14185 => "01101010", 14188 => "01110101", 14194 => "11101001", 14195 => "01100110", 14196 => "00101101", 14197 => "01110111", 14198 => "00001011", 14200 => "01100001", 14202 => "10111010", 14203 => "11100011", 14204 => "01011101", 14209 => "01110000", 14211 => "01011011", 14212 => "10001110", 14214 => "10000000", 14216 => "00000111", 14217 => "11111001", 14218 => "00000110", 14221 => "00111000", 14222 => "10011001", 14223 => "10111011", 14224 => "10010110", 14225 => "11000001", 14227 => "10101000", 14230 => "10011000", 14233 => "01010000", 14234 => "10010111", 14238 => "01100001", 14239 => "10000000", 14241 => "11101110", 14242 => "11101010", 14243 => "10111100", 14244 => "11110010", 14245 => "00010001", 14247 => "10010000", 14250 => "10000100", 14251 => "01001110", 14256 => "11001001", 14257 => "10011101", 14258 => "10000011", 14261 => "00001110", 14262 => "11001011", 14263 => "01010010", 14265 => "10111100", 14267 => "00001011", 14268 => "10101110", 14269 => "00010101", 14270 => "10100101", 14271 => "10111110", 14276 => "11110011", 14279 => "11111010", 14280 => "00000011", 14281 => "11001010", 14283 => "10011000", 14284 => "10111111", 14285 => "10011011", 14286 => "01011110", 14290 => "01010010", 14291 => "00100111", 14299 => "11101101", 14300 => "11101110", 14301 => "01001001", 14303 => "10011000", 14304 => "00001101", 14306 => "01000001", 14307 => "00010110", 14311 => "11101101", 14314 => "10100011", 14316 => "00110110", 14319 => "11101011", 14320 => "00010001", 14322 => "00100010", 14324 => "00010011", 14326 => "11111000", 14327 => "11100101", 14329 => "10010100", 14330 => "11000000", 14334 => "01000110", 14335 => "01101011", 14340 => "11101100", 14341 => "10100100", 14349 => "00001001", 14351 => "01100011", 14354 => "10100111", 14356 => "00101111", 14357 => "10001111", 14358 => "10011010", 14360 => "01011100", 14362 => "11111110", 14364 => "01100101", 14365 => "10100000", 14367 => "00010101", 14368 => "10100100", 14371 => "11011001", 14372 => "10101111", 14373 => "01010100", 14374 => "10110111", 14377 => "01111101", 14379 => "00001111", 14380 => "10011011", 14381 => "11100111", 14382 => "11111010", 14383 => "10000110", 14384 => "11011110", 14388 => "01110000", 14392 => "11000111", 14394 => "01111110", 14397 => "11010100", 14402 => "00000101", 14403 => "01010000", 14405 => "00111110", 14408 => "10110100", 14409 => "00011111", 14412 => "01011111", 14413 => "11101100", 14414 => "00011101", 14416 => "00001011", 14417 => "10011110", 14418 => "11011101", 14424 => "10000010", 14429 => "00010010", 14431 => "00111100", 14434 => "01010110", 14435 => "01001101", 14436 => "11011100", 14440 => "00000100", 14441 => "10010111", 14442 => "01010100", 14446 => "10010000", 14447 => "10001111", 14448 => "01101100", 14449 => "00001101", 14450 => "00001011", 14451 => "10100111", 14454 => "10010010", 14459 => "00001001", 14463 => "00000001", 14466 => "10010010", 14468 => "11001101", 14472 => "00001110", 14473 => "00100001", 14474 => "00100011", 14475 => "00100010", 14477 => "01111101", 14479 => "11101111", 14485 => "11110001", 14486 => "11110010", 14488 => "10100101", 14489 => "11010011", 14491 => "00011011", 14498 => "01010010", 14499 => "10100010", 14505 => "01101010", 14507 => "10000000", 14508 => "01111110", 14509 => "01001000", 14510 => "10010000", 14512 => "10010010", 14513 => "10101010", 14516 => "01110110", 14518 => "11001100", 14519 => "10011110", 14521 => "10100110", 14527 => "10100010", 14529 => "11010110", 14530 => "00010011", 14533 => "10000100", 14536 => "10010010", 14538 => "01101001", 14544 => "01010001", 14545 => "11100001", 14548 => "10110010", 14550 => "10111000", 14551 => "10110001", 14555 => "10010001", 14560 => "01001101", 14562 => "11101111", 14563 => "11111000", 14568 => "10011010", 14569 => "00101010", 14572 => "00010101", 14574 => "11001100", 14579 => "10000000", 14581 => "11110101", 14584 => "00101011", 14586 => "00010001", 14589 => "00100110", 14590 => "00000001", 14591 => "01111011", 14594 => "01010010", 14597 => "10110000", 14598 => "01111011", 14599 => "10100100", 14604 => "11011100", 14605 => "11011000", 14607 => "00100000", 14609 => "00101100", 14615 => "10111100", 14617 => "11100110", 14618 => "01010001", 14619 => "01100011", 14622 => "00011111", 14624 => "01011001", 14625 => "01010000", 14626 => "00111111", 14627 => "10011010", 14631 => "11111110", 14633 => "00001111", 14634 => "11000011", 14639 => "11000000", 14640 => "01011101", 14645 => "00001110", 14646 => "10001111", 14647 => "11111101", 14648 => "11000001", 14649 => "01111101", 14650 => "11110101", 14652 => "10100111", 14656 => "00101011", 14657 => "00110111", 14658 => "11100110", 14660 => "00100011", 14662 => "11100101", 14665 => "01000000", 14666 => "00000001", 14667 => "10000010", 14669 => "11110100", 14670 => "11000111", 14672 => "11110111", 14674 => "11010110", 14675 => "10011111", 14676 => "01111111", 14677 => "01011010", 14678 => "11001010", 14680 => "00011001", 14682 => "11101001", 14684 => "10001011", 14687 => "10101100", 14688 => "00010100", 14690 => "00010110", 14693 => "11011111", 14694 => "00111001", 14696 => "10111111", 14697 => "10101010", 14699 => "00001111", 14701 => "00111011", 14708 => "00111001", 14709 => "11100101", 14711 => "11110110", 14717 => "00001000", 14719 => "01110111", 14722 => "10101110", 14724 => "10001010", 14726 => "01100000", 14727 => "10011011", 14728 => "10000000", 14729 => "11100010", 14730 => "10100101", 14731 => "10110001", 14732 => "01011111", 14733 => "01010111", 14735 => "11110110", 14736 => "11111100", 14738 => "00101111", 14741 => "10110010", 14742 => "01111100", 14744 => "10111011", 14745 => "01001000", 14749 => "01100100", 14750 => "01111000", 14752 => "11010000", 14755 => "01111011", 14756 => "11101000", 14762 => "11000010", 14763 => "10110111", 14765 => "11101001", 14768 => "01100101", 14775 => "10000011", 14777 => "00011010", 14781 => "10111011", 14782 => "00000111", 14784 => "00100100", 14785 => "10010011", 14786 => "00110101", 14789 => "11011100", 14791 => "01111101", 14797 => "00010000", 14801 => "11111100", 14804 => "00110101", 14805 => "00001110", 14808 => "01000101", 14811 => "01110111", 14812 => "01111100", 14813 => "01001111", 14820 => "11111110", 14821 => "11110001", 14823 => "11110110", 14825 => "01100100", 14826 => "11001100", 14827 => "01110011", 14828 => "11010001", 14829 => "01111111", 14830 => "11001101", 14833 => "01011100", 14834 => "00111011", 14835 => "00100100", 14840 => "10100001", 14841 => "11111001", 14843 => "11110110", 14844 => "11111010", 14845 => "00011010", 14847 => "10110000", 14848 => "10110000", 14851 => "10001001", 14854 => "01110001", 14855 => "10011111", 14857 => "00101110", 14858 => "11101110", 14862 => "11010100", 14863 => "10011111", 14866 => "01000000", 14869 => "11000000", 14872 => "01011010", 14873 => "01100000", 14874 => "11001111", 14878 => "00010011", 14879 => "10101110", 14880 => "01000100", 14881 => "10011000", 14882 => "11100111", 14886 => "10001111", 14887 => "01011110", 14889 => "11011101", 14890 => "01111110", 14892 => "10001110", 14895 => "01101010", 14897 => "01010001", 14899 => "01101100", 14900 => "01101101", 14902 => "11010010", 14903 => "00101000", 14905 => "00111011", 14906 => "00010100", 14914 => "10100110", 14916 => "10111000", 14919 => "01010100", 14920 => "10111011", 14921 => "10001001", 14924 => "10011110", 14926 => "10100001", 14930 => "01000010", 14938 => "00011001", 14941 => "11001011", 14944 => "11000111", 14946 => "10001101", 14947 => "00000010", 14948 => "00000010", 14949 => "10100110", 14950 => "11000011", 14951 => "10010110", 14952 => "01100001", 14954 => "10111110", 14959 => "10100110", 14968 => "00101000", 14969 => "10010001", 14971 => "01001111", 14976 => "00010000", 14977 => "00011010", 14979 => "11001001", 14980 => "10011100", 14989 => "00010011", 14990 => "01011100", 14991 => "00111010", 14992 => "01101101", 14993 => "01001111", 14997 => "01111010", 14999 => "11100100", 15000 => "11000100", 15001 => "10111010", 15003 => "01110100", 15006 => "10010100", 15008 => "00000001", 15009 => "10100100", 15010 => "10011010", 15011 => "01011010", 15012 => "00000100", 15014 => "00101101", 15015 => "10101000", 15016 => "10110110", 15019 => "10100101", 15021 => "01000110", 15022 => "11001110", 15023 => "10001000", 15028 => "01110000", 15030 => "11001001", 15031 => "10110011", 15032 => "10101000", 15033 => "11010011", 15034 => "00011000", 15035 => "00011101", 15037 => "01000001", 15038 => "00010101", 15039 => "11111101", 15041 => "10010011", 15042 => "10100101", 15044 => "00010011", 15045 => "00000101", 15048 => "01011000", 15049 => "11110010", 15052 => "00111100", 15055 => "11101101", 15056 => "10100011", 15059 => "01101010", 15061 => "10100111", 15064 => "00000011", 15070 => "11110010", 15071 => "10011000", 15076 => "10100011", 15080 => "00010000", 15081 => "01001011", 15083 => "10000101", 15085 => "11001001", 15086 => "00100101", 15087 => "10001110", 15088 => "00100111", 15090 => "01001100", 15094 => "10011011", 15097 => "10001000", 15098 => "00100111", 15100 => "11110100", 15103 => "01100110", 15106 => "00100111", 15108 => "10111111", 15110 => "11110100", 15112 => "11001010", 15113 => "11111110", 15114 => "00010101", 15123 => "11100001", 15124 => "00111000", 15125 => "11111000", 15126 => "11101001", 15129 => "00100001", 15130 => "10101101", 15132 => "01100111", 15133 => "01000001", 15138 => "01011001", 15140 => "00110111", 15141 => "10011111", 15142 => "00011000", 15143 => "00110000", 15144 => "01001101", 15145 => "00110110", 15147 => "01101111", 15149 => "10101110", 15150 => "00010010", 15153 => "10001001", 15157 => "01100011", 15160 => "10100001", 15161 => "11100001", 15163 => "11001010", 15168 => "11101110", 15169 => "01100000", 15173 => "10110001", 15174 => "11000111", 15175 => "01000010", 15176 => "00000011", 15178 => "10001011", 15184 => "01000111", 15185 => "00111101", 15186 => "11001100", 15192 => "10101110", 15195 => "00111101", 15196 => "01110010", 15198 => "00111100", 15205 => "01000000", 15206 => "10111111", 15208 => "11000110", 15212 => "01110111", 15213 => "11111111", 15216 => "11000000", 15218 => "11001001", 15220 => "00111101", 15221 => "01111001", 15222 => "00011101", 15223 => "00000001", 15224 => "01011011", 15225 => "01001111", 15228 => "11011101", 15229 => "10001000", 15230 => "11101010", 15233 => "00010111", 15235 => "00001111", 15236 => "11000010", 15238 => "00101111", 15240 => "00100011", 15242 => "00110100", 15246 => "01010110", 15247 => "00100100", 15248 => "10010000", 15252 => "11111101", 15255 => "00001000", 15256 => "00111110", 15257 => "10110100", 15258 => "00101110", 15260 => "10100000", 15261 => "01111011", 15262 => "01001010", 15264 => "10111100", 15265 => "01101100", 15267 => "10001011", 15268 => "01100101", 15269 => "00101011", 15273 => "00100010", 15276 => "10001000", 15277 => "11010111", 15281 => "11111111", 15282 => "11000101", 15284 => "00010011", 15285 => "01001001", 15286 => "01101111", 15287 => "01001011", 15288 => "10010001", 15291 => "01100101", 15293 => "00001011", 15296 => "11110001", 15297 => "00100000", 15298 => "11000001", 15299 => "01100110", 15301 => "01100001", 15302 => "10111010", 15307 => "01011101", 15308 => "10111100", 15312 => "01011111", 15314 => "11000001", 15315 => "11111111", 15316 => "10100101", 15320 => "11100101", 15322 => "00100101", 15325 => "10011011", 15327 => "10101110", 15328 => "00000111", 15329 => "01110100", 15332 => "00110111", 15333 => "00010000", 15336 => "10100010", 15339 => "01100000", 15344 => "00011110", 15345 => "10001001", 15349 => "00100110", 15354 => "00111110", 15355 => "01111111", 15357 => "11010000", 15358 => "01100101", 15360 => "10111100", 15361 => "01100000", 15364 => "00011101", 15365 => "00111101", 15368 => "11011111", 15371 => "01000111", 15372 => "10010011", 15375 => "11000001", 15379 => "11110010", 15384 => "00000111", 15385 => "00101111", 15390 => "11110100", 15392 => "01110111", 15394 => "11101100", 15395 => "10110001", 15396 => "00101100", 15397 => "01000011", 15399 => "11101110", 15404 => "11000100", 15405 => "10101101", 15406 => "00111010", 15407 => "01011110", 15408 => "10001000", 15410 => "11000001", 15413 => "11100101", 15416 => "00001110", 15417 => "01111110", 15421 => "01010111", 15426 => "01110101", 15428 => "10011011", 15429 => "10110101", 15433 => "10001101", 15434 => "00001110", 15437 => "00111100", 15438 => "11001001", 15439 => "11111110", 15443 => "01110011", 15448 => "11001110", 15450 => "01001011", 15451 => "01000101", 15452 => "01110001", 15453 => "11101100", 15454 => "11101100", 15456 => "00101001", 15459 => "01011010", 15461 => "00010010", 15462 => "01100110", 15464 => "01011111", 15465 => "01101100", 15466 => "10100010", 15467 => "01110101", 15468 => "11101110", 15474 => "11110000", 15475 => "01101001", 15476 => "01110100", 15477 => "00010001", 15478 => "00010000", 15480 => "10001101", 15482 => "11110110", 15485 => "01011111", 15486 => "01000110", 15491 => "01111001", 15492 => "11101010", 15494 => "00000101", 15497 => "10010100", 15498 => "01011111", 15499 => "00111100", 15503 => "00111101", 15504 => "10001111", 15506 => "11100111", 15507 => "11100010", 15508 => "00011010", 15509 => "01101101", 15511 => "10100111", 15514 => "11011111", 15515 => "10001011", 15518 => "10011010", 15519 => "01001001", 15520 => "11000110", 15521 => "01100000", 15524 => "00110110", 15525 => "11100000", 15530 => "00100001", 15531 => "11110011", 15532 => "10000110", 15536 => "10110010", 15539 => "01101001", 15540 => "10011101", 15541 => "10011100", 15545 => "01001100", 15546 => "01100000", 15548 => "00001100", 15551 => "10011010", 15552 => "01000010", 15553 => "01010010", 15557 => "00010110", 15558 => "00010100", 15563 => "10011101", 15564 => "11100000", 15565 => "10011000", 15566 => "01010010", 15568 => "10000100", 15569 => "01010010", 15572 => "10011010", 15576 => "11001101", 15578 => "10011000", 15580 => "11011011", 15581 => "11110100", 15582 => "10001001", 15584 => "01010011", 15586 => "00100000", 15587 => "01100111", 15592 => "01100110", 15593 => "11010101", 15594 => "11010101", 15600 => "11001000", 15605 => "00111110", 15607 => "10010011", 15608 => "11110100", 15613 => "11101110", 15614 => "01011001", 15616 => "10011100", 15617 => "10100001", 15618 => "01100011", 15619 => "10011001", 15621 => "00111010", 15622 => "01110000", 15624 => "11001000", 15626 => "11110111", 15627 => "10000110", 15629 => "01110100", 15630 => "00011110", 15631 => "11110111", 15632 => "11100111", 15635 => "00011101", 15641 => "01010011", 15642 => "01011010", 15643 => "11111001", 15647 => "01111011", 15650 => "11111001", 15652 => "11110110", 15654 => "11111101", 15655 => "11000001", 15656 => "11101011", 15660 => "10111001", 15663 => "00010101", 15665 => "10000111", 15666 => "10000111", 15667 => "00001100", 15669 => "10001111", 15670 => "01110001", 15674 => "11101111", 15676 => "11000100", 15677 => "00011000", 15684 => "10011110", 15685 => "01010110", 15686 => "10101011", 15687 => "11110011", 15689 => "01100111", 15690 => "11110100", 15691 => "11011111", 15692 => "11001000", 15698 => "00111100", 15700 => "11000111", 15701 => "01101101", 15702 => "11110101", 15703 => "01000100", 15705 => "01010011", 15706 => "00101110", 15707 => "11000111", 15715 => "00111110", 15716 => "10001000", 15717 => "01110110", 15718 => "11111100", 15719 => "11100110", 15720 => "01111101", 15721 => "11101101", 15722 => "00100100", 15724 => "10010011", 15725 => "11010100", 15726 => "11010011", 15727 => "10110011", 15728 => "11011001", 15734 => "11110011", 15741 => "00100011", 15742 => "11111000", 15745 => "11100010", 15746 => "11101011", 15747 => "01011001", 15748 => "00010101", 15749 => "00011100", 15751 => "11101100", 15756 => "11001010", 15759 => "11111000", 15760 => "01001010", 15761 => "11001110", 15766 => "01111110", 15767 => "10011000", 15768 => "11100110", 15770 => "11010100", 15777 => "01001010", 15778 => "11010101", 15780 => "01011100", 15781 => "01011010", 15783 => "10000101", 15784 => "11110011", 15789 => "00111010", 15790 => "11011010", 15793 => "00000010", 15794 => "00011100", 15797 => "10000010", 15798 => "11010001", 15805 => "00001010", 15806 => "00010101", 15807 => "11000000", 15810 => "11110111", 15811 => "10110010", 15815 => "10000011", 15816 => "00101001", 15817 => "11111110", 15819 => "11100110", 15821 => "00101100", 15823 => "10000000", 15825 => "01111100", 15827 => "10100111", 15828 => "10111001", 15830 => "11100010", 15831 => "10001100", 15834 => "00111100", 15835 => "10101000", 15838 => "01110001", 15843 => "00011001", 15844 => "00010010", 15847 => "01010111", 15850 => "10111100", 15851 => "10000101", 15852 => "01111100", 15855 => "10101101", 15856 => "00100010", 15858 => "11110101", 15865 => "01001010", 15867 => "10111110", 15870 => "10000101", 15871 => "10111000", 15872 => "10000111", 15875 => "01011110", 15879 => "01100001", 15881 => "00001110", 15883 => "11011101", 15888 => "01111011", 15890 => "10111000", 15891 => "00111100", 15894 => "00111000", 15896 => "00011000", 15898 => "00000011", 15899 => "01100011", 15900 => "01101010", 15902 => "00000110", 15906 => "11011111", 15907 => "11000001", 15909 => "10000001", 15910 => "00000010", 15913 => "00001000", 15916 => "00010101", 15918 => "01110110", 15920 => "10101000", 15922 => "11001111", 15925 => "01011100", 15926 => "11010011", 15927 => "10011100", 15929 => "11111101", 15931 => "10000111", 15932 => "11100110", 15933 => "00100011", 15934 => "00110010", 15936 => "01000110", 15938 => "00111111", 15940 => "01100001", 15942 => "00101011", 15955 => "01010100", 15959 => "00111000", 15961 => "10001011", 15965 => "00011011", 15966 => "11010011", 15967 => "11111010", 15968 => "11001110", 15970 => "00110011", 15972 => "10001010", 15973 => "11101010", 15974 => "10101100", 15975 => "10111000", 15976 => "00111011", 15977 => "00101001", 15978 => "01101010", 15981 => "00110000", 15982 => "11010101", 15985 => "10000101", 15986 => "00100001", 15988 => "00011010", 15991 => "01010011", 15993 => "00011110", 15994 => "11000111", 15995 => "00000011", 15997 => "10100011", 15999 => "10001010", 16003 => "11110010", 16004 => "01101111", 16006 => "11100110", 16011 => "00001011", 16015 => "01010100", 16017 => "00001101", 16018 => "11100011", 16020 => "11101000", 16022 => "00101001", 16024 => "01100010", 16027 => "10001100", 16028 => "10111010", 16035 => "01001100", 16039 => "11011100", 16041 => "11111010", 16045 => "10011101", 16047 => "01011010", 16049 => "11101100", 16050 => "10001011", 16053 => "00111001", 16056 => "10101001", 16061 => "01110000", 16062 => "00001010", 16064 => "10100100", 16072 => "00100111", 16073 => "00001111", 16075 => "01101111", 16076 => "00111001", 16077 => "11101011", 16083 => "10111000", 16085 => "11001010", 16087 => "01111101", 16089 => "01001101", 16091 => "00001100", 16094 => "11100101", 16095 => "11100010", 16097 => "11110110", 16098 => "11001111", 16099 => "10110000", 16100 => "10100010", 16102 => "11001010", 16103 => "01111110", 16106 => "11001001", 16107 => "00001111", 16109 => "10101101", 16110 => "10010011", 16111 => "00110111", 16112 => "00000100", 16114 => "01010101", 16115 => "11001010", 16119 => "00010111", 16120 => "10110000", 16126 => "01011000", 16135 => "01000011", 16137 => "10010001", 16142 => "11011111", 16145 => "01010111", 16146 => "01111010", 16147 => "10111110", 16148 => "00100111", 16149 => "10110100", 16151 => "11011011", 16152 => "11110111", 16153 => "00100011", 16154 => "10111100", 16155 => "11110100", 16156 => "11111011", 16157 => "11100001", 16162 => "11001000", 16163 => "10010100", 16166 => "11000001", 16167 => "01111101", 16171 => "11000000", 16172 => "10111010", 16175 => "11011111", 16178 => "00010001", 16179 => "01000011", 16180 => "00110000", 16181 => "01001010", 16182 => "00010000", 16184 => "10010111", 16185 => "10000010", 16186 => "01000011", 16187 => "00000011", 16189 => "10101001", 16193 => "00000011", 16197 => "10011001", 16199 => "11011010", 16200 => "11111101", 16201 => "01001100", 16202 => "00000001", 16205 => "11111101", 16206 => "10011101", 16207 => "00000001", 16209 => "00101111", 16210 => "11001101", 16214 => "01000101", 16215 => "00101000", 16216 => "11101100", 16218 => "10111011", 16219 => "10011100", 16220 => "10001110", 16222 => "10001011", 16223 => "00101110", 16224 => "10010010", 16226 => "11000010", 16227 => "11011000", 16228 => "11100110", 16234 => "01010000", 16236 => "00011100", 16237 => "10011100", 16241 => "10000101", 16245 => "10110011", 16246 => "10011001", 16247 => "10000101", 16248 => "00001011", 16250 => "01010000", 16251 => "11100011", 16256 => "01001101", 16258 => "01111101", 16261 => "11001100", 16262 => "11100010", 16263 => "10000100", 16268 => "11101010", 16269 => "00011010", 16272 => "10110101", 16274 => "01100100", 16276 => "10101111", 16282 => "01100111", 16283 => "01011100", 16285 => "01001000", 16287 => "01000100", 16291 => "01111111", 16293 => "01010110", 16296 => "01100010", 16298 => "01000111", 16305 => "01101100", 16306 => "11000010", 16307 => "01110101", 16310 => "10000000", 16316 => "11010010", 16317 => "10000111", 16320 => "01101101", 16322 => "11010111", 16324 => "00101101", 16326 => "11010001", 16331 => "10110001", 16334 => "10101100", 16336 => "01111011", 16338 => "01100110", 16344 => "11010111", 16346 => "11100010", 16347 => "01010101", 16348 => "11010100", 16349 => "01001100", 16350 => "10101100", 16352 => "10010110", 16356 => "00100111", 16357 => "10101000", 16358 => "11010101", 16360 => "11001111", 16361 => "01111110", 16364 => "01111001", 16365 => "10001101", 16374 => "01000111", 16375 => "10000110", 16377 => "01110011", 16379 => "00110101", 16381 => "00011110", 16382 => "01101010", 16386 => "11101110", 16389 => "11011001", 16392 => "10101011", 16394 => "00000101", 16396 => "00111011", 16398 => "00101110", 16399 => "11000110", 16407 => "10111001", 16408 => "01011100", 16409 => "11010110", 16412 => "11000001", 16413 => "00110110", 16415 => "11001011", 16416 => "10010000", 16420 => "00110011", 16421 => "11110110", 16423 => "00100001", 16425 => "11010011", 16429 => "10011111", 16436 => "10101000", 16439 => "00100000", 16440 => "00110100", 16442 => "11000101", 16443 => "11100011", 16445 => "01110011", 16446 => "10000100", 16447 => "01110110", 16448 => "10100100", 16449 => "10010110", 16452 => "01111011", 16453 => "00010010", 16455 => "01001110", 16456 => "11110101", 16457 => "11110000", 16458 => "01111011", 16459 => "11110100", 16460 => "11000011", 16462 => "11110011", 16463 => "01010111", 16464 => "00001010", 16465 => "11101010", 16467 => "01011010", 16468 => "11101111", 16470 => "11011100", 16473 => "01010011", 16475 => "00111010", 16476 => "10000000", 16479 => "11100011", 16480 => "00100110", 16483 => "00101111", 16486 => "11011100", 16489 => "01010101", 16491 => "11001001", 16494 => "00110111", 16500 => "01001110", 16502 => "01101101", 16503 => "00010110", 16505 => "01110011", 16508 => "01000100", 16515 => "01111011", 16516 => "11101111", 16518 => "10011111", 16520 => "00010001", 16522 => "11101111", 16523 => "11100001", 16525 => "10100010", 16529 => "10101100", 16531 => "10100001", 16532 => "10000101", 16534 => "10011010", 16535 => "10011001", 16537 => "11111110", 16542 => "11100000", 16543 => "01011111", 16544 => "00001111", 16545 => "11101100", 16546 => "00010010", 16547 => "10011100", 16553 => "00010111", 16554 => "01001000", 16557 => "01110010", 16560 => "01100111", 16566 => "01110000", 16567 => "00100001", 16569 => "11011111", 16575 => "00010001", 16576 => "11110101", 16579 => "00101001", 16582 => "00111001", 16584 => "11101100", 16585 => "01000001", 16586 => "10110011", 16587 => "00001011", 16590 => "00110110", 16593 => "01101100", 16594 => "00001110", 16598 => "11101000", 16599 => "01100010", 16601 => "11010100", 16603 => "11011111", 16605 => "11010110", 16608 => "10000101", 16609 => "10101110", 16611 => "10010101", 16612 => "10001001", 16616 => "10001111", 16617 => "10001010", 16618 => "11101000", 16619 => "11110011", 16621 => "10101100", 16624 => "01111110", 16627 => "01001011", 16629 => "11111000", 16630 => "10011000", 16631 => "01011000", 16633 => "10101101", 16634 => "01000111", 16636 => "00100110", 16637 => "01011010", 16638 => "01011010", 16639 => "10011111", 16641 => "00111001", 16642 => "00110111", 16643 => "11101000", 16644 => "00010000", 16645 => "11100111", 16648 => "00001011", 16650 => "00111110", 16652 => "11101111", 16653 => "00101010", 16655 => "11011001", 16658 => "11011111", 16662 => "01010001", 16663 => "10001101", 16666 => "00111110", 16668 => "00001101", 16669 => "11001001", 16672 => "11100101", 16673 => "00100111", 16676 => "10000011", 16679 => "11111011", 16680 => "00110101", 16681 => "10010000", 16682 => "10100101", 16683 => "00001001", 16684 => "01110010", 16685 => "10100110", 16687 => "11111001", 16688 => "11101111", 16690 => "00001101", 16692 => "10100100", 16694 => "11100001", 16697 => "01000010", 16699 => "01010001", 16700 => "10101011", 16701 => "01001001", 16702 => "00011101", 16704 => "00100010", 16705 => "01010111", 16707 => "10011001", 16709 => "10010101", 16710 => "01100000", 16711 => "00000110", 16713 => "11000010", 16714 => "01011010", 16718 => "11010101", 16719 => "10100010", 16720 => "01110010", 16723 => "11110000", 16724 => "11111010", 16725 => "01001001", 16727 => "00000100", 16729 => "10100010", 16730 => "11101010", 16733 => "11001001", 16735 => "10000100", 16736 => "10101110", 16737 => "00010010", 16738 => "11000001", 16739 => "11111001", 16740 => "10011111", 16743 => "01100001", 16744 => "01111000", 16745 => "10010101", 16746 => "10010101", 16749 => "11011000", 16751 => "11011110", 16752 => "00100111", 16754 => "00010100", 16756 => "11101000", 16758 => "10110110", 16759 => "01101100", 16761 => "00100101", 16764 => "01001000", 16765 => "11000000", 16769 => "11111111", 16770 => "01001010", 16777 => "00011101", 16778 => "01011011", 16779 => "11011111", 16781 => "10000000", 16782 => "00001001", 16783 => "11000010", 16784 => "11011000", 16795 => "10000010", 16796 => "10000010", 16800 => "01011000", 16801 => "00000100", 16804 => "10111100", 16806 => "10000010", 16812 => "00110111", 16821 => "10110101", 16822 => "11000110", 16823 => "11111011", 16824 => "01110100", 16827 => "11101010", 16832 => "00101001", 16833 => "11000101", 16836 => "00101001", 16839 => "11010011", 16840 => "00010000", 16841 => "00100111", 16844 => "11011100", 16846 => "01101111", 16847 => "00010001", 16848 => "00010011", 16849 => "10110001", 16853 => "00100010", 16854 => "00111001", 16858 => "00110001", 16859 => "10111101", 16860 => "11001010", 16861 => "11110010", 16862 => "10110111", 16863 => "00110110", 16865 => "00001110", 16868 => "00001010", 16869 => "11000011", 16871 => "01101000", 16873 => "01110011", 16876 => "11010101", 16883 => "11000000", 16884 => "11011110", 16888 => "00010100", 16891 => "11001100", 16892 => "01001000", 16893 => "11001011", 16894 => "01001110", 16895 => "11001111", 16896 => "00101001", 16904 => "01001000", 16905 => "01010101", 16908 => "00111101", 16910 => "01001111", 16912 => "10111011", 16914 => "01001100", 16917 => "10001000", 16920 => "11000111", 16924 => "11100110", 16925 => "00111101", 16928 => "00111000", 16929 => "00000110", 16930 => "00100101", 16931 => "11001101", 16933 => "10111001", 16934 => "11001100", 16936 => "10110011", 16938 => "10111001", 16940 => "11000011", 16943 => "01100100", 16945 => "01000111", 16946 => "01010011", 16948 => "11111110", 16949 => "01001010", 16953 => "01001101", 16954 => "00010001", 16956 => "11001001", 16958 => "01101110", 16962 => "01010011", 16963 => "01101011", 16964 => "01100110", 16968 => "11101101", 16970 => "01101011", 16971 => "00100100", 16973 => "01000100", 16974 => "10101101", 16978 => "10011101", 16979 => "10011101", 16980 => "01010011", 16981 => "11101010", 16984 => "11000000", 16985 => "01010000", 16986 => "11101101", 16987 => "00110111", 16992 => "01101101", 16993 => "01101100", 16994 => "01111010", 16996 => "00000111", 16998 => "00011001", 17000 => "00110110", 17003 => "00010001", 17006 => "11101100", 17007 => "10011101", 17008 => "10101101", 17009 => "11001010", 17011 => "00110000", 17013 => "10101111", 17014 => "01001010", 17015 => "10101000", 17016 => "10001100", 17019 => "11011000", 17020 => "00100100", 17022 => "00111001", 17023 => "10100111", 17025 => "00011000", 17029 => "00101000", 17030 => "01100001", 17031 => "10011111", 17035 => "00101101", 17040 => "01101100", 17041 => "10110100", 17043 => "10111001", 17044 => "01111111", 17045 => "00001011", 17046 => "10101110", 17047 => "11101111", 17049 => "10011011", 17050 => "01110010", 17054 => "10111000", 17055 => "10110011", 17060 => "01101111", 17062 => "10111001", 17064 => "10101001", 17065 => "01001010", 17066 => "11101100", 17068 => "10011110", 17069 => "11000010", 17070 => "11011111", 17071 => "11110011", 17073 => "10110001", 17077 => "10010010", 17083 => "01001111", 17086 => "10101001", 17087 => "00101010", 17089 => "00111111", 17091 => "11110111", 17092 => "11011000", 17094 => "11001111", 17097 => "00111011", 17099 => "10001010", 17100 => "01101010", 17101 => "10111101", 17102 => "10100100", 17105 => "11110100", 17106 => "01111011", 17107 => "01011110", 17112 => "01100111", 17115 => "00001110", 17117 => "10011000", 17120 => "01011001", 17121 => "01111101", 17122 => "00100010", 17127 => "00101001", 17129 => "10110010", 17134 => "01001010", 17135 => "00101001", 17144 => "10000101", 17148 => "11001011", 17150 => "11110100", 17151 => "10011000", 17152 => "10110111", 17153 => "00000101", 17154 => "00001010", 17157 => "11010111", 17161 => "00010101", 17163 => "01101001", 17170 => "10001110", 17171 => "00001010", 17172 => "11100000", 17175 => "01011011", 17176 => "11110010", 17178 => "11011110", 17179 => "00111011", 17181 => "11100110", 17187 => "11010101", 17188 => "10111100", 17189 => "01100110", 17191 => "11101100", 17192 => "00011100", 17193 => "10100100", 17194 => "11010101", 17197 => "01010111", 17198 => "00110010", 17201 => "00000011", 17202 => "00101111", 17205 => "11001110", 17206 => "01110010", 17207 => "11110100", 17210 => "01100111", 17215 => "10011000", 17223 => "00011111", 17224 => "00010010", 17225 => "00011001", 17226 => "00000111", 17227 => "00001110", 17229 => "01101011", 17234 => "00001100", 17235 => "00100011", 17236 => "11010011", 17237 => "10110111", 17240 => "10111100", 17242 => "10110000", 17243 => "01010101", 17244 => "11111010", 17245 => "11100001", 17246 => "00010100", 17250 => "10010010", 17252 => "00101001", 17255 => "00010000", 17256 => "11110001", 17259 => "01011000", 17262 => "11011111", 17264 => "10011001", 17267 => "01110100", 17268 => "10010010", 17269 => "10011011", 17270 => "11111001", 17271 => "01001000", 17273 => "11111110", 17277 => "00111111", 17280 => "11011011", 17283 => "01100010", 17285 => "01101000", 17288 => "10010010", 17289 => "11100110", 17290 => "01101111", 17291 => "01001100", 17293 => "01010110", 17294 => "11101111", 17295 => "01000000", 17296 => "00110111", 17300 => "10110111", 17303 => "01111011", 17305 => "10110001", 17306 => "01000101", 17309 => "00111000", 17311 => "10000010", 17313 => "10000101", 17314 => "11111000", 17316 => "10100101", 17320 => "00010110", 17322 => "10111110", 17323 => "11100010", 17325 => "11110100", 17327 => "01000101", 17329 => "01011101", 17330 => "01110100", 17331 => "10100011", 17335 => "01011111", 17336 => "00001111", 17347 => "10110010", 17348 => "00111100", 17349 => "01101101", 17350 => "10011110", 17352 => "11100101", 17357 => "11111100", 17359 => "10100011", 17363 => "01110111", 17364 => "11110001", 17369 => "10110110", 17371 => "11010011", 17373 => "11101001", 17375 => "00011000", 17376 => "10110011", 17377 => "11100000", 17378 => "11001101", 17382 => "00011111", 17383 => "10011111", 17384 => "10011110", 17389 => "00110010", 17390 => "01010011", 17391 => "11000100", 17393 => "10100110", 17395 => "11110100", 17396 => "01011001", 17397 => "01100001", 17400 => "01110011", 17402 => "10100001", 17405 => "00000011", 17407 => "10100100", 17409 => "01010000", 17410 => "10000010", 17411 => "10111111", 17412 => "10100110", 17414 => "10000110", 17420 => "10000110", 17422 => "00001110", 17425 => "11000100", 17428 => "11100110", 17429 => "11101010", 17434 => "10111010", 17440 => "10111010", 17441 => "00010000", 17443 => "00011000", 17444 => "01111000", 17445 => "10010001", 17446 => "11100000", 17448 => "11000101", 17450 => "01100010", 17451 => "11111010", 17456 => "11101100", 17459 => "10101001", 17460 => "11100110", 17463 => "11010111", 17464 => "10011000", 17465 => "11010010", 17466 => "01100010", 17472 => "01010011", 17473 => "10110000", 17476 => "10100010", 17477 => "11011111", 17481 => "01101000", 17483 => "10001101", 17484 => "00010101", 17485 => "00000110", 17488 => "00001011", 17490 => "01111101", 17492 => "11010101", 17493 => "10110100", 17494 => "11001100", 17496 => "01111001", 17497 => "11101110", 17498 => "00111001", 17499 => "10110110", 17502 => "11000010", 17503 => "11000101", 17504 => "10011110", 17507 => "10110110", 17512 => "01100001", 17514 => "01111001", 17516 => "00100111", 17517 => "01011101", 17519 => "10011111", 17523 => "11101010", 17524 => "10001110", 17525 => "10000010", 17526 => "00010011", 17528 => "00100111", 17530 => "10011111", 17531 => "00110000", 17535 => "01111100", 17537 => "00111000", 17540 => "01010000", 17541 => "00101111", 17542 => "11011100", 17544 => "10000101", 17547 => "11001011", 17554 => "00010100", 17557 => "11011010", 17558 => "00101001", 17559 => "10101000", 17563 => "00000111", 17564 => "10101000", 17571 => "00011110", 17572 => "10001100", 17573 => "11011010", 17575 => "10100111", 17577 => "00111011", 17579 => "11000000", 17582 => "10111010", 17587 => "00000010", 17588 => "11001101", 17589 => "01011111", 17591 => "11111111", 17593 => "01000101", 17594 => "01011010", 17595 => "10000101", 17597 => "01111000", 17600 => "11111101", 17601 => "11011000", 17603 => "00011111", 17607 => "11010110", 17608 => "10111000", 17612 => "01110000", 17613 => "11000100", 17616 => "00101101", 17618 => "00000011", 17619 => "00100000", 17620 => "10000001", 17622 => "01001100", 17626 => "01100001", 17627 => "00101000", 17629 => "10110110", 17630 => "01111000", 17632 => "00111000", 17633 => "01010111", 17635 => "11110011", 17636 => "00010110", 17637 => "10011011", 17641 => "10100110", 17646 => "01111110", 17647 => "11100111", 17648 => "01101100", 17652 => "11101111", 17653 => "11110000", 17656 => "00110110", 17657 => "10010001", 17659 => "10101110", 17660 => "10111011", 17661 => "01110010", 17662 => "11011110", 17665 => "10010111", 17666 => "10000101", 17671 => "10111010", 17672 => "10011011", 17678 => "11010000", 17680 => "00101100", 17681 => "01100001", 17682 => "00010100", 17683 => "10111100", 17686 => "10100101", 17687 => "00101000", 17689 => "00010011", 17690 => "01010000", 17693 => "00111100", 17694 => "11111011", 17696 => "10101010", 17699 => "00011101", 17701 => "01110000", 17704 => "00010100", 17706 => "01100101", 17707 => "10000100", 17712 => "11001000", 17713 => "10110001", 17715 => "11011010", 17716 => "10011001", 17718 => "01000010", 17719 => "00010101", 17722 => "01100001", 17724 => "01000000", 17726 => "00101111", 17727 => "11101110", 17728 => "10110101", 17730 => "01101001", 17731 => "00100110", 17733 => "10000000", 17734 => "10101100", 17737 => "11000111", 17741 => "10101100", 17742 => "11000000", 17743 => "01111001", 17747 => "11110111", 17750 => "10111111", 17751 => "11111010", 17754 => "01101010", 17756 => "00100100", 17757 => "00100000", 17759 => "11110000", 17761 => "11111001", 17762 => "11111101", 17767 => "01000001", 17773 => "11000010", 17774 => "10010000", 17775 => "10100000", 17776 => "00000110", 17781 => "11001000", 17782 => "10101011", 17785 => "11111101", 17787 => "01011111", 17789 => "11100000", 17791 => "10011011", 17792 => "01110100", 17794 => "10010100", 17795 => "11110101", 17796 => "11111110", 17798 => "10010011", 17799 => "01100001", 17800 => "01110010", 17803 => "10110000", 17804 => "11000101", 17806 => "11111001", 17811 => "11100001", 17812 => "10011001", 17813 => "00010101", 17815 => "10011100", 17817 => "10011101", 17820 => "00100000", 17823 => "10100100", 17824 => "00111100", 17825 => "01001110", 17830 => "11011000", 17838 => "00110111", 17839 => "10001011", 17841 => "11001100", 17842 => "00110111", 17844 => "10001010", 17845 => "10111010", 17846 => "10001010", 17847 => "11101111", 17848 => "11110011", 17849 => "01010101", 17850 => "01101011", 17851 => "01110111", 17853 => "00011111", 17854 => "10011000", 17855 => "01001100", 17856 => "01001000", 17858 => "11010110", 17860 => "00001100", 17862 => "10110010", 17864 => "00111111", 17866 => "01111111", 17867 => "11111101", 17868 => "11011001", 17870 => "11011110", 17873 => "11101001", 17875 => "00001001", 17878 => "00001101", 17879 => "00011010", 17882 => "01000110", 17884 => "01111100", 17887 => "11110101", 17889 => "00111110", 17891 => "11001101", 17893 => "01001010", 17894 => "00110101", 17895 => "00011111", 17898 => "00010100", 17903 => "01111110", 17904 => "00000001", 17906 => "00101110", 17907 => "11001110", 17908 => "11010010", 17909 => "01000010", 17910 => "00000011", 17914 => "11101000", 17916 => "01110101", 17917 => "10110101", 17920 => "10110010", 17924 => "00000100", 17925 => "00101000", 17928 => "01100101", 17929 => "10101010", 17930 => "10000001", 17932 => "10011000", 17934 => "01011011", 17936 => "10011011", 17938 => "10101001", 17939 => "11010011", 17941 => "01011110", 17942 => "01101010", 17946 => "01100110", 17950 => "11111001", 17951 => "00011101", 17954 => "01001111", 17955 => "01001011", 17960 => "10111100", 17962 => "10011000", 17966 => "01000100", 17967 => "00111010", 17968 => "11101110", 17969 => "01011000", 17970 => "11011110", 17974 => "01101011", 17975 => "00110001", 17979 => "10001101", 17981 => "00011011", 17982 => "01110011", 17983 => "10000101", 17984 => "00100100", 17986 => "10111110", 17987 => "11000110", 17988 => "01111000", 17989 => "11110001", 17990 => "10001101", 17991 => "11011100", 17993 => "11100000", 17994 => "10100010", 17997 => "00011110", 17998 => "00010111", 18000 => "01101111", 18001 => "01001111", 18002 => "00111110", 18004 => "10100111", 18005 => "10000110", 18009 => "00110110", 18011 => "10010010", 18012 => "00011010", 18014 => "00101001", 18015 => "01000010", 18019 => "10001101", 18023 => "11011110", 18025 => "11011000", 18026 => "01010110", 18027 => "10100001", 18032 => "00010000", 18033 => "10001100", 18035 => "11011011", 18037 => "00101101", 18038 => "10100000", 18039 => "00111111", 18040 => "10100101", 18042 => "01000101", 18050 => "10100000", 18051 => "11101000", 18052 => "11011011", 18053 => "00001010", 18058 => "01001110", 18059 => "00011010", 18061 => "10100100", 18066 => "00010001", 18070 => "10010101", 18071 => "01001100", 18077 => "10101100", 18078 => "01001111", 18082 => "11110011", 18083 => "11111101", 18084 => "01011110", 18085 => "10111001", 18086 => "00011100", 18089 => "10000010", 18092 => "11001110", 18094 => "10100110", 18096 => "01101000", 18099 => "10110010", 18103 => "00110011", 18105 => "10100111", 18108 => "00011000", 18109 => "00010111", 18114 => "10000101", 18115 => "01100111", 18118 => "10001000", 18121 => "11100110", 18125 => "10010101", 18126 => "00010110", 18127 => "10011101", 18130 => "01001011", 18133 => "11010101", 18134 => "10001101", 18135 => "10111100", 18137 => "10001110", 18138 => "00111111", 18141 => "11101011", 18142 => "11011110", 18143 => "11011111", 18147 => "01111000", 18149 => "11111111", 18152 => "11010010", 18153 => "00011010", 18157 => "10011010", 18159 => "10011010", 18160 => "10110011", 18162 => "01110010", 18163 => "00101010", 18165 => "01110001", 18173 => "01101111", 18174 => "11110101", 18175 => "10000000", 18176 => "11000111", 18178 => "10111111", 18179 => "10010010", 18180 => "00111001", 18182 => "00100101", 18184 => "00110011", 18187 => "00111110", 18191 => "11010100", 18195 => "11011111", 18199 => "11100001", 18200 => "01011000", 18201 => "01100110", 18203 => "10000001", 18206 => "00001101", 18207 => "01101100", 18208 => "11001011", 18209 => "11101111", 18213 => "01000111", 18214 => "00100010", 18215 => "00001010", 18219 => "11011000", 18221 => "00100110", 18224 => "01110000", 18225 => "01100011", 18227 => "00110001", 18229 => "00001011", 18231 => "10101100", 18239 => "01000001", 18240 => "10110011", 18241 => "01100110", 18244 => "01111101", 18245 => "00000001", 18247 => "00000010", 18248 => "01001011", 18250 => "00111010", 18253 => "00110001", 18257 => "10101110", 18259 => "00000101", 18261 => "10011111", 18262 => "01101101", 18263 => "01001110", 18264 => "11001110", 18265 => "01100101", 18267 => "01100111", 18269 => "01001011", 18271 => "01101100", 18272 => "11101000", 18275 => "10011101", 18276 => "00000011", 18278 => "01001010", 18280 => "01100111", 18282 => "10101100", 18283 => "01110111", 18284 => "01111111", 18286 => "11100100", 18290 => "00101010", 18293 => "00101101", 18294 => "00010100", 18299 => "00101001", 18301 => "10001010", 18303 => "11110001", 18304 => "01000110", 18305 => "10010001", 18309 => "00110101", 18313 => "01011000", 18314 => "11111010", 18315 => "01111010", 18317 => "00001000", 18318 => "10010101", 18320 => "10000110", 18322 => "10000000", 18324 => "10101011", 18326 => "00100000", 18327 => "01110101", 18329 => "01111000", 18331 => "10111000", 18332 => "11001001", 18334 => "00001111", 18336 => "01101001", 18339 => "01001100", 18342 => "01110110", 18346 => "01100000", 18347 => "00101110", 18348 => "00000101", 18350 => "11111011", 18352 => "01001011", 18353 => "01110000", 18354 => "01111101", 18356 => "00001101", 18357 => "11010101", 18358 => "10101000", 18361 => "01000110", 18362 => "01000101", 18364 => "00110110", 18365 => "10111001", 18369 => "10101101", 18370 => "10100101", 18374 => "01011001", 18375 => "11010111", 18376 => "10000100", 18381 => "11011110", 18382 => "01101111", 18386 => "01010011", 18389 => "11101001", 18391 => "00001101", 18395 => "11010011", 18398 => "01010001", 18399 => "00010100", 18400 => "11000111", 18401 => "10010001", 18407 => "00001111", 18409 => "00110001", 18411 => "11100001", 18412 => "10100010", 18414 => "10011100", 18416 => "01011011", 18422 => "10011011", 18425 => "10111000", 18426 => "11100011", 18427 => "00001101", 18431 => "11001010", 18437 => "00011111", 18439 => "01011001", 18441 => "11101101", 18443 => "00001011", 18446 => "00111000", 18448 => "10000000", 18451 => "10001101", 18452 => "11101101", 18453 => "10111110", 18454 => "10101011", 18457 => "11011100", 18461 => "00001001", 18464 => "00011001", 18466 => "00101010", 18467 => "01110101", 18468 => "01101111", 18469 => "10000101", 18473 => "11011001", 18474 => "00011100", 18483 => "01101011", 18484 => "01111001", 18486 => "00100100", 18488 => "00110011", 18494 => "01101101", 18496 => "10101100", 18497 => "11110110", 18500 => "00111100", 18501 => "10010100", 18503 => "11110110", 18505 => "00111010", 18506 => "00001011", 18507 => "11111110", 18510 => "10010100", 18511 => "10011001", 18513 => "00001111", 18514 => "01111101", 18516 => "11000111", 18517 => "10111100", 18518 => "11000110", 18519 => "11010011", 18520 => "00100100", 18524 => "01111001", 18525 => "00000110", 18526 => "01000001", 18527 => "00100011", 18529 => "01111101", 18530 => "10001011", 18531 => "10001010", 18536 => "01010010", 18537 => "00010111", 18538 => "01010001", 18539 => "11001001", 18545 => "01000000", 18546 => "11111110", 18548 => "11010000", 18550 => "00111110", 18551 => "10001111", 18553 => "10101010", 18557 => "11111000", 18558 => "00010000", 18563 => "01111111", 18565 => "01110001", 18567 => "10000010", 18568 => "10111111", 18569 => "10111111", 18570 => "11010010", 18572 => "11011111", 18576 => "11001001", 18581 => "00101010", 18583 => "11010010", 18584 => "01011110", 18585 => "10111100", 18587 => "11110110", 18592 => "11010010", 18593 => "10100111", 18598 => "01110110", 18600 => "11011110", 18602 => "11010001", 18604 => "01110001", 18605 => "10110111", 18606 => "00111110", 18608 => "01010100", 18609 => "11000011", 18610 => "11011011", 18613 => "00111011", 18619 => "10111010", 18622 => "01100101", 18624 => "10000111", 18625 => "01011100", 18626 => "00101110", 18627 => "01100101", 18628 => "10011011", 18631 => "11101001", 18636 => "01001011", 18637 => "00111011", 18644 => "11000000", 18648 => "11100100", 18649 => "00101000", 18651 => "00001110", 18653 => "01111001", 18655 => "10001000", 18656 => "00101011", 18658 => "10110110", 18659 => "00110100", 18661 => "11110100", 18666 => "01010010", 18669 => "01000100", 18670 => "01010110", 18671 => "00111111", 18677 => "10111110", 18678 => "00101001", 18679 => "00011110", 18682 => "10011000", 18683 => "01011001", 18685 => "10010110", 18686 => "00111000", 18689 => "00001001", 18691 => "00101111", 18692 => "10110110", 18697 => "10110110", 18699 => "10110010", 18701 => "10011110", 18703 => "01101110", 18705 => "00101001", 18706 => "00001101", 18708 => "00111010", 18710 => "01110000", 18711 => "01001110", 18713 => "10000000", 18717 => "01011101", 18718 => "10010101", 18719 => "10000001", 18720 => "11001000", 18721 => "11111011", 18723 => "01001001", 18724 => "01110111", 18727 => "11100101", 18730 => "01010010", 18731 => "11010000", 18732 => "01100001", 18734 => "10000001", 18735 => "00101000", 18737 => "11011011", 18738 => "01111100", 18739 => "01011111", 18740 => "01101011", 18742 => "00001110", 18746 => "00000001", 18747 => "00101111", 18750 => "11111001", 18751 => "01001111", 18755 => "11111000", 18762 => "11000001", 18765 => "11101001", 18769 => "01010110", 18772 => "11011110", 18774 => "10110110", 18775 => "00111001", 18776 => "00101100", 18779 => "10101011", 18780 => "01101011", 18783 => "11001110", 18786 => "00111001", 18787 => "11011111", 18788 => "01100010", 18791 => "00001101", 18794 => "01011001", 18795 => "01011010", 18796 => "10011010", 18797 => "01001001", 18798 => "01011100", 18800 => "11101111", 18802 => "00111000", 18805 => "00010000", 18806 => "01111000", 18808 => "01000101", 18809 => "11101011", 18815 => "11111001", 18817 => "01001100", 18819 => "10001110", 18820 => "01101001", 18821 => "10000000", 18822 => "00000110", 18823 => "00101101", 18825 => "11001000", 18826 => "01011111", 18828 => "01100010", 18830 => "01101101", 18831 => "10100011", 18832 => "00010101", 18835 => "01000101", 18836 => "01111011", 18837 => "10100100", 18844 => "11000010", 18846 => "11011001", 18847 => "11111101", 18848 => "10000100", 18849 => "11101010", 18850 => "10101111", 18852 => "11101001", 18854 => "11000100", 18855 => "01110011", 18857 => "10111010", 18858 => "10011011", 18862 => "01000110", 18865 => "11101011", 18867 => "01001001", 18870 => "00100100", 18871 => "00010100", 18872 => "00100101", 18874 => "11000001", 18880 => "01110111", 18883 => "11011000", 18885 => "11000010", 18888 => "10000100", 18891 => "01010111", 18893 => "00001011", 18894 => "01001101", 18895 => "11010011", 18897 => "00100010", 18898 => "01000011", 18899 => "10111101", 18900 => "00011101", 18903 => "11010100", 18904 => "11010001", 18905 => "00010110", 18907 => "11010011", 18908 => "11110100", 18911 => "10001101", 18917 => "11110001", 18918 => "10100100", 18919 => "11110111", 18922 => "00101111", 18923 => "01001110", 18926 => "11001101", 18927 => "00101100", 18933 => "11001000", 18934 => "10100111", 18937 => "10111111", 18939 => "11111110", 18941 => "11001100", 18942 => "11001110", 18946 => "11100101", 18948 => "00001101", 18950 => "10100111", 18952 => "11100000", 18953 => "10011000", 18954 => "00110100", 18956 => "11110000", 18960 => "10101101", 18961 => "10100111", 18962 => "01011010", 18964 => "11011110", 18966 => "01001110", 18967 => "01000110", 18968 => "11011110", 18970 => "01001101", 18971 => "01111101", 18972 => "01101101", 18975 => "00001001", 18977 => "01010100", 18978 => "11001100", 18980 => "01000001", 18981 => "11101001", 18983 => "11000110", 18984 => "10001011", 18987 => "10100100", 18988 => "10101110", 18989 => "11000000", 18990 => "11111010", 18994 => "10001001", 18996 => "11000001", 18999 => "01000001", 19001 => "11110010", 19002 => "11001101", 19003 => "11011000", 19006 => "11001111", 19007 => "00011000", 19011 => "10001010", 19014 => "00011011", 19019 => "10110110", 19020 => "11000000", 19021 => "10100000", 19023 => "11001111", 19026 => "11011011", 19027 => "01110000", 19028 => "01110001", 19034 => "00010110", 19035 => "11010110", 19036 => "01001001", 19037 => "01101000", 19038 => "00100001", 19041 => "10101011", 19042 => "00010110", 19043 => "10010011", 19047 => "10100100", 19048 => "11101100", 19056 => "00001111", 19063 => "01110101", 19064 => "10011110", 19068 => "10001000", 19069 => "00000111", 19070 => "01100000", 19072 => "11100101", 19073 => "00101101", 19074 => "10001010", 19076 => "01110110", 19077 => "01111010", 19078 => "11010110", 19079 => "00010011", 19081 => "01101010", 19083 => "00010100", 19084 => "01001100", 19086 => "10111100", 19087 => "00000110", 19089 => "00111111", 19090 => "00101010", 19091 => "01110100", 19092 => "11011100", 19095 => "01110101", 19096 => "01010111", 19097 => "01011101", 19098 => "10011100", 19101 => "11100101", 19102 => "10110101", 19103 => "01111001", 19105 => "11111010", 19109 => "01001011", 19111 => "01000010", 19113 => "01111110", 19116 => "11010010", 19117 => "11000111", 19118 => "00100110", 19121 => "11010010", 19122 => "00100010", 19125 => "10001101", 19126 => "10110000", 19127 => "01010110", 19128 => "10001010", 19129 => "10000001", 19130 => "00000001", 19131 => "10011001", 19134 => "10001011", 19135 => "00010010", 19137 => "11100100", 19138 => "11100101", 19139 => "10111100", 19141 => "10000110", 19142 => "10110010", 19144 => "10110110", 19147 => "10011001", 19150 => "11110111", 19151 => "10111010", 19154 => "00110101", 19155 => "10100010", 19162 => "00000010", 19163 => "11110011", 19165 => "10100110", 19166 => "00001111", 19168 => "00101100", 19171 => "00000110", 19172 => "10100110", 19173 => "10101100", 19175 => "00111000", 19178 => "10110110", 19179 => "10111111", 19181 => "11000011", 19182 => "00001110", 19183 => "10111111", 19184 => "01001000", 19185 => "00011101", 19187 => "01110011", 19195 => "01001101", 19196 => "11010011", 19197 => "01000000", 19199 => "00100101", 19202 => "01001101", 19203 => "11001100", 19208 => "10000001", 19209 => "00100100", 19211 => "10011010", 19214 => "01111000", 19219 => "01100000", 19220 => "01111010", 19223 => "11111010", 19224 => "11111110", 19225 => "00111110", 19228 => "11000000", 19229 => "10101011", 19230 => "00010010", 19236 => "11111101", 19240 => "10001101", 19242 => "11010110", 19244 => "10010100", 19246 => "10110000", 19249 => "10001110", 19250 => "01001110", 19251 => "11110011", 19252 => "00110100", 19257 => "00110110", 19263 => "00101000", 19265 => "11110011", 19268 => "01001100", 19272 => "01011111", 19274 => "10011111", 19277 => "11011010", 19278 => "00111100", 19279 => "01011010", 19280 => "01011101", 19281 => "00001110", 19283 => "11000001", 19285 => "01010110", 19286 => "01001110", 19288 => "10100011", 19290 => "10011000", 19303 => "01111100", 19304 => "11100000", 19305 => "10001111", 19306 => "11110111", 19308 => "10111110", 19309 => "01101111", 19312 => "00010001", 19316 => "01110010", 19318 => "10110101", 19320 => "11000111", 19321 => "01111101", 19322 => "10010101", 19323 => "01111010", 19330 => "01101001", 19333 => "01111110", 19334 => "10011000", 19335 => "01100000", 19336 => "01001110", 19338 => "10001100", 19339 => "11000110", 19340 => "10101000", 19344 => "11010011", 19345 => "01111010", 19346 => "00001100", 19349 => "11110100", 19354 => "11111011", 19357 => "10010011", 19359 => "00010011", 19362 => "01001001", 19364 => "00111001", 19365 => "11001000", 19367 => "10011111", 19368 => "01110111", 19372 => "01011111", 19374 => "00101010", 19375 => "01010100", 19379 => "10110000", 19380 => "10110111", 19381 => "11000101", 19382 => "00111000", 19384 => "10000001", 19385 => "10101110", 19386 => "10110010", 19388 => "10010111", 19389 => "00000010", 19391 => "11100001", 19392 => "00110010", 19396 => "01010011", 19397 => "00001001", 19398 => "01101011", 19399 => "10100111", 19403 => "01011101", 19407 => "01100101", 19409 => "11100111", 19410 => "11110110", 19413 => "01011110", 19414 => "00001001", 19417 => "11100001", 19418 => "10111001", 19419 => "10000110", 19421 => "10101101", 19422 => "00011111", 19423 => "00100001", 19424 => "00100111", 19425 => "01100000", 19427 => "10000100", 19428 => "00001001", 19429 => "01100111", 19431 => "11110011", 19432 => "00001100", 19433 => "10010010", 19434 => "01011011", 19435 => "10011111", 19436 => "01010010", 19438 => "11111100", 19441 => "00000100", 19442 => "10000110", 19446 => "01101101", 19448 => "00010010", 19449 => "01111110", 19450 => "10001010", 19455 => "11101010", 19457 => "01100100", 19458 => "00101001", 19461 => "10011101", 19462 => "11110111", 19464 => "11111000", 19465 => "11011100", 19466 => "01001001", 19469 => "11111011", 19470 => "11001010", 19471 => "10011011", 19476 => "10101000", 19477 => "10000000", 19480 => "11110010", 19481 => "01110001", 19483 => "00011011", 19485 => "00100111", 19489 => "11011011", 19491 => "11100110", 19495 => "00001011", 19496 => "11011010", 19498 => "00110110", 19499 => "01000010", 19500 => "10010000", 19503 => "11110010", 19506 => "11001010", 19508 => "01000001", 19510 => "10110001", 19511 => "11000010", 19513 => "10111110", 19515 => "00100010", 19517 => "01000001", 19518 => "00100010", 19519 => "01110011", 19521 => "10100011", 19524 => "00001000", 19525 => "00001110", 19526 => "10000011", 19528 => "10100010", 19530 => "11101000", 19531 => "10011000", 19532 => "00010100", 19534 => "00110010", 19535 => "11110101", 19537 => "01001101", 19540 => "11100101", 19541 => "00000100", 19543 => "00111000", 19545 => "00000011", 19547 => "01000011", 19549 => "01110001", 19552 => "01101100", 19554 => "00001000", 19561 => "10001101", 19562 => "11101010", 19563 => "10101000", 19564 => "10111000", 19565 => "00010010", 19566 => "01100011", 19570 => "10001111", 19575 => "10111100", 19577 => "00010100", 19579 => "00010011", 19580 => "11010111", 19582 => "10110100", 19586 => "11010110", 19587 => "00111110", 19588 => "01011101", 19594 => "10110010", 19595 => "00000111", 19596 => "11111100", 19599 => "01001110", 19600 => "00101110", 19601 => "00000100", 19602 => "10100100", 19603 => "11110000", 19606 => "01000011", 19612 => "01111101", 19613 => "11000100", 19614 => "01111001", 19615 => "10001101", 19616 => "10000000", 19620 => "10111100", 19625 => "01101000", 19627 => "01100010", 19629 => "10001101", 19630 => "00000100", 19631 => "01101110", 19633 => "10010101", 19634 => "01001001", 19635 => "10111100", 19638 => "00101100", 19639 => "11001000", 19640 => "11001101", 19642 => "01110111", 19643 => "00100000", 19645 => "01001011", 19650 => "10001001", 19651 => "10110111", 19652 => "00011111", 19653 => "01001100", 19655 => "10100101", 19656 => "01011100", 19657 => "00101000", 19658 => "01000001", 19661 => "11000000", 19662 => "11110101", 19663 => "11000110", 19665 => "00011101", 19667 => "10100101", 19668 => "11010011", 19669 => "10001100", 19670 => "10000011", 19671 => "00010101", 19674 => "10101010", 19677 => "01000100", 19687 => "11111100", 19689 => "00011111", 19692 => "10100110", 19693 => "10011001", 19695 => "01110000", 19697 => "11111001", 19700 => "10110110", 19701 => "10100001", 19711 => "00100111", 19712 => "10111011", 19717 => "01110101", 19721 => "00111011", 19722 => "10000110", 19727 => "01010000", 19728 => "00100011", 19729 => "10101011", 19732 => "10101001", 19735 => "11110010", 19736 => "00101001", 19739 => "00100001", 19740 => "01001101", 19741 => "10010101", 19743 => "01101110", 19744 => "11110100", 19747 => "11010111", 19748 => "11011010", 19749 => "10001010", 19750 => "01100111", 19752 => "01111010", 19755 => "11010001", 19756 => "11000000", 19758 => "10101111", 19760 => "01010100", 19761 => "00111011", 19763 => "00000011", 19764 => "01111001", 19765 => "00110101", 19766 => "11001111", 19767 => "10010111", 19771 => "00011101", 19777 => "01111000", 19780 => "01111011", 19781 => "10011100", 19783 => "00110011", 19788 => "10000011", 19791 => "11000010", 19792 => "01111100", 19795 => "01010001", 19796 => "01001101", 19799 => "11010001", 19800 => "00110001", 19802 => "00100100", 19803 => "00110000", 19804 => "00101100", 19808 => "10111111", 19810 => "00100001", 19811 => "00111111", 19812 => "00000110", 19816 => "11111010", 19817 => "00011101", 19822 => "00101110", 19825 => "00111000", 19829 => "01100010", 19833 => "11010000", 19834 => "11111010", 19836 => "00000001", 19840 => "00010010", 19841 => "00101001", 19846 => "10111010", 19850 => "11111100", 19851 => "01111101", 19854 => "10110011", 19855 => "00001001", 19856 => "11000100", 19857 => "11101010", 19859 => "00010101", 19861 => "10101001", 19864 => "10111101", 19865 => "10101110", 19866 => "11110000", 19872 => "00011101", 19874 => "01001001", 19876 => "11100000", 19878 => "11011001", 19883 => "01111110", 19886 => "11010110", 19888 => "10101010", 19889 => "11001111", 19890 => "00001110", 19891 => "01101000", 19896 => "10010010", 19897 => "10001101", 19899 => "10111011", 19901 => "11000000", 19902 => "10011101", 19903 => "01001100", 19905 => "11100010", 19909 => "00000011", 19912 => "00010001", 19917 => "11000010", 19920 => "01010111", 19922 => "10100111", 19925 => "11010101", 19928 => "10001110", 19932 => "00111011", 19934 => "10000001", 19935 => "00100100", 19937 => "10100110", 19938 => "00110001", 19939 => "11111000", 19941 => "00110001", 19943 => "10000001", 19947 => "11110001", 19948 => "01110011", 19949 => "00001000", 19950 => "00111011", 19952 => "11110000", 19955 => "00100111", 19956 => "11101111", 19960 => "10001110", 19962 => "00110011", 19968 => "01010000", 19969 => "11110011", 19970 => "11110001", 19971 => "10001101", 19972 => "10001101", 19973 => "11110101", 19974 => "01001110", 19976 => "11001101", 19977 => "01111000", 19982 => "01001100", 19987 => "10011010", 19988 => "11010000", 19990 => "11000010", 19994 => "11000100", 19995 => "01011111", 20000 => "00101100", 20003 => "00011110", 20004 => "01110010", 20006 => "10100111", 20008 => "00101111", 20009 => "11111001", 20010 => "10100101", 20014 => "10101100", 20015 => "00110110", 20017 => "00011001", 20019 => "11001011", 20020 => "11110111", 20024 => "10011101", 20026 => "10101010", 20029 => "00001011", 20030 => "11001101", 20031 => "01011000", 20032 => "10101101", 20033 => "00111010", 20036 => "10010101", 20039 => "11011001", 20041 => "01101101", 20047 => "01011110", 20048 => "11001011", 20049 => "10011011", 20050 => "11110001", 20052 => "00010000", 20056 => "01010011", 20058 => "10011011", 20059 => "10101110", 20061 => "11110001", 20062 => "10000100", 20068 => "01101100", 20070 => "11111100", 20072 => "00010011", 20073 => "11011111", 20074 => "11000000", 20075 => "00111101", 20077 => "01010010", 20079 => "00000101", 20084 => "11111000", 20086 => "01011100", 20087 => "01010000", 20090 => "10110101", 20093 => "10010101", 20096 => "10110101", 20099 => "10101001", 20100 => "00101101", 20102 => "10111011", 20104 => "01000110", 20105 => "11001001", 20109 => "10001110", 20110 => "11001101", 20115 => "00100010", 20116 => "01011001", 20117 => "00101000", 20119 => "01000011", 20121 => "10010111", 20123 => "00101011", 20126 => "11110111", 20127 => "00111110", 20128 => "10100001", 20130 => "11011101", 20132 => "10011100", 20134 => "00001000", 20135 => "01011111", 20138 => "11010011", 20143 => "11011001", 20144 => "00100110", 20145 => "00010001", 20146 => "00011110", 20147 => "00011100", 20148 => "00101010", 20149 => "01011111", 20150 => "01010001", 20152 => "10110000", 20153 => "10010000", 20155 => "01001110", 20156 => "00100001", 20158 => "01011011", 20159 => "10101111", 20160 => "01000000", 20162 => "10101100", 20163 => "10001101", 20164 => "01110100", 20165 => "01001001", 20167 => "11010101", 20171 => "01010111", 20175 => "10111000", 20177 => "10000000", 20178 => "10100000", 20179 => "01100100", 20181 => "01110100", 20191 => "11100001", 20192 => "01000101", 20193 => "00011111", 20194 => "00010111", 20195 => "00001000", 20197 => "10001000", 20201 => "11000110", 20204 => "10100001", 20207 => "00101011", 20208 => "00111000", 20211 => "00001011", 20215 => "00001100", 20218 => "10001101", 20219 => "00001100", 20220 => "01011000", 20221 => "10100100", 20225 => "00010010", 20229 => "00111110", 20233 => "00101010", 20244 => "01001010", 20247 => "10100110", 20248 => "00000011", 20249 => "11100110", 20251 => "01101100", 20252 => "01011110", 20253 => "11110010", 20257 => "00010001", 20258 => "10101110", 20263 => "00110100", 20264 => "01110000", 20266 => "01100010", 20267 => "01100110", 20268 => "00001101", 20270 => "01000000", 20271 => "11100010", 20272 => "10010110", 20273 => "00111011", 20276 => "01100110", 20277 => "00111111", 20278 => "11011101", 20282 => "01110100", 20283 => "10011001", 20285 => "11110100", 20287 => "00111101", 20288 => "00011101", 20289 => "11011010", 20292 => "11101000", 20296 => "01111011", 20299 => "10100101", 20302 => "01010000", 20303 => "10010101", 20304 => "11001010", 20312 => "10110110", 20313 => "10101010", 20314 => "11100000", 20315 => "10000011", 20316 => "10001001", 20317 => "00010010", 20320 => "01000011", 20323 => "01111011", 20324 => "01110011", 20325 => "10010001", 20326 => "01111110", 20328 => "01100001", 20331 => "11100101", 20332 => "11110011", 20333 => "10101111", 20334 => "10111100", 20335 => "11001000", 20337 => "10000100", 20340 => "01010100", 20342 => "10101000", 20343 => "10000110", 20346 => "00011010", 20349 => "11100101", 20350 => "10011110", 20353 => "00101100", 20354 => "00111010", 20355 => "00100001", 20356 => "11100010", 20358 => "00111001", 20361 => "10100100", 20366 => "11000101", 20367 => "01100000", 20369 => "00110100", 20371 => "10001010", 20372 => "10111111", 20374 => "10101101", 20376 => "00001010", 20378 => "00111011", 20382 => "01000100", 20384 => "10111101", 20385 => "01011111", 20386 => "10111100", 20387 => "00110100", 20389 => "00000010", 20392 => "00100110", 20395 => "01011000", 20398 => "11100001", 20399 => "10111011", 20402 => "10111110", 20403 => "11000010", 20404 => "00100100", 20407 => "10101110", 20408 => "00110111", 20412 => "10001101", 20415 => "01010110", 20416 => "11100111", 20420 => "10111101", 20422 => "11001101", 20423 => "10010111", 20424 => "11000111", 20429 => "10001111", 20430 => "00110111", 20431 => "01011001", 20432 => "11000001", 20433 => "11000101", 20434 => "10101000", 20435 => "11101100", 20440 => "01101001", 20444 => "00010000", 20449 => "01000001", 20450 => "10110010", 20455 => "11110010", 20460 => "01110101", 20461 => "01111011", 20465 => "11111000", 20467 => "01001011", 20468 => "10111010", 20469 => "10101001", 20471 => "01010011", 20472 => "10011100", 20473 => "10111101", 20474 => "01000111", 20478 => "11100000", 20480 => "10101101", 20481 => "01011011", 20483 => "10011010", 20484 => "11000110", 20488 => "10010001", 20489 => "00001001", 20490 => "10000010", 20492 => "10101010", 20493 => "10110000", 20495 => "11110000", 20496 => "00010100", 20498 => "01000111", 20499 => "01111001", 20500 => "01111010", 20503 => "11101101", 20506 => "11001110", 20507 => "10111101", 20508 => "00011110", 20509 => "11100010", 20510 => "10111010", 20513 => "01011010", 20514 => "11110101", 20515 => "10111000", 20516 => "10111110", 20522 => "10111010", 20525 => "00101001", 20527 => "11111011", 20529 => "01000101", 20530 => "11001110", 20535 => "01011011", 20538 => "10111101", 20539 => "11011110", 20540 => "10101110", 20542 => "00100011", 20544 => "11011001", 20545 => "11101001", 20546 => "11100001", 20549 => "11001111", 20550 => "01110010", 20551 => "00110110", 20552 => "10101101", 20554 => "10111011", 20555 => "00100001", 20556 => "01010011", 20563 => "00101001", 20564 => "11011001", 20565 => "11111000", 20568 => "10100011", 20572 => "01010110", 20574 => "01100010", 20580 => "10111101", 20581 => "11011011", 20585 => "00100001", 20586 => "01111001", 20587 => "00001011", 20590 => "01010100", 20591 => "11001100", 20592 => "11001100", 20594 => "10000100", 20595 => "11011111", 20596 => "11011100", 20597 => "10100111", 20598 => "11010000", 20602 => "10101000", 20603 => "00011100", 20608 => "01011100", 20611 => "11001000", 20612 => "10111110", 20613 => "11010100", 20622 => "10110011", 20623 => "01111000", 20625 => "10111010", 20626 => "00100011", 20630 => "00110101", 20636 => "11000111", 20641 => "11110011", 20643 => "11101011", 20645 => "10110101", 20646 => "10100101", 20648 => "00111110", 20650 => "10010101", 20652 => "11100010", 20654 => "10110010", 20656 => "10100000", 20657 => "11000110", 20658 => "00110001", 20661 => "10111110", 20662 => "10001111", 20663 => "01010111", 20664 => "10001011", 20666 => "01010000", 20670 => "11100111", 20673 => "01011001", 20675 => "11110101", 20676 => "10101110", 20680 => "00000001", 20686 => "01000001", 20688 => "01011001", 20695 => "00101111", 20697 => "11101100", 20698 => "10100000", 20702 => "00110110", 20705 => "01011111", 20707 => "01000010", 20708 => "11000101", 20710 => "11100111", 20711 => "00000101", 20714 => "10000000", 20717 => "11101011", 20718 => "10110101", 20719 => "11010000", 20720 => "11011000", 20721 => "00011111", 20722 => "00101010", 20723 => "11011010", 20724 => "10000011", 20726 => "00000011", 20727 => "00001100", 20729 => "10101010", 20732 => "00001011", 20733 => "11111000", 20736 => "00100001", 20739 => "10111000", 20740 => "11101101", 20741 => "00000011", 20744 => "11111001", 20746 => "01001101", 20753 => "10111001", 20754 => "01100010", 20755 => "10010010", 20764 => "10001001", 20765 => "01101010", 20768 => "11010001", 20769 => "11110100", 20770 => "10000111", 20773 => "00010001", 20775 => "11100111", 20778 => "00010011", 20779 => "11111101", 20781 => "00101101", 20782 => "01001111", 20784 => "11001110", 20787 => "00111010", 20790 => "11101101", 20791 => "00100101", 20792 => "00010100", 20795 => "00110101", 20796 => "01101010", 20799 => "01010000", 20804 => "11100010", 20805 => "01010101", 20807 => "00111101", 20811 => "11110000", 20814 => "10010110", 20815 => "11101010", 20817 => "10111101", 20819 => "00100000", 20820 => "01111001", 20823 => "01101010", 20827 => "10001111", 20828 => "10000110", 20831 => "11000001", 20836 => "10001011", 20840 => "01000000", 20845 => "11110100", 20846 => "01011011", 20847 => "00000001", 20848 => "00001011", 20850 => "11101000", 20852 => "00111000", 20857 => "10100111", 20858 => "01100000", 20859 => "01010010", 20861 => "01000000", 20867 => "11111101", 20868 => "10101100", 20873 => "10110000", 20877 => "00101010", 20882 => "10010100", 20885 => "11010100", 20887 => "00010100", 20888 => "10110111", 20891 => "01010011", 20892 => "10001010", 20895 => "11001010", 20897 => "01010001", 20898 => "01011010", 20899 => "10011111", 20902 => "11000001", 20904 => "11011011", 20905 => "00001010", 20906 => "10010110", 20907 => "00010011", 20909 => "00001001", 20911 => "01000010", 20912 => "01011001", 20913 => "00110011", 20914 => "10000000", 20915 => "10110111", 20919 => "11101000", 20921 => "00101011", 20922 => "01011010", 20926 => "00110011", 20934 => "01101011", 20935 => "00011001", 20939 => "11111000", 20941 => "10110101", 20942 => "01000111", 20943 => "00010110", 20944 => "10111000", 20946 => "01010110", 20947 => "10100110", 20948 => "01000011", 20949 => "10000101", 20950 => "10001100", 20953 => "00100010", 20954 => "01010001", 20958 => "00011000", 20960 => "00101110", 20962 => "01100101", 20963 => "10010001", 20964 => "00011000", 20965 => "11000100", 20969 => "10000010", 20972 => "01100010", 20973 => "01001011", 20974 => "00110000", 20977 => "00010000", 20978 => "10011101", 20979 => "11011100", 20981 => "00100101", 20985 => "00110011", 20988 => "11000001", 20989 => "11101010", 20990 => "11110010", 20991 => "00011101", 20992 => "01001100", 20993 => "01110110", 20995 => "10111110", 20996 => "00000111", 20998 => "00000100", 21000 => "11011001", 21001 => "00011000", 21002 => "00001110", 21003 => "00110110", 21005 => "10111000", 21008 => "01011000", 21009 => "00001100", 21010 => "11100001", 21018 => "10110010", 21020 => "10110011", 21021 => "01000001", 21022 => "11111011", 21024 => "01011110", 21025 => "01100010", 21027 => "00001000", 21028 => "00010101", 21029 => "11101010", 21030 => "01001010", 21034 => "11110000", 21035 => "01111101", 21036 => "01110110", 21038 => "11000111", 21044 => "00000100", 21046 => "00011001", 21047 => "00010011", 21049 => "11110111", 21050 => "01001110", 21055 => "11101000", 21056 => "10011011", 21057 => "00100110", 21059 => "11000100", 21062 => "11011111", 21065 => "10101100", 21066 => "11110011", 21071 => "11101101", 21072 => "10101110", 21075 => "10001001", 21076 => "00100111", 21077 => "11101100", 21080 => "01110111", 21086 => "11010111", 21088 => "00000011", 21090 => "00111111", 21091 => "10010000", 21094 => "00100111", 21095 => "11110000", 21096 => "01110100", 21098 => "11000101", 21101 => "11010010", 21103 => "00001011", 21104 => "11110100", 21105 => "11110000", 21107 => "01111010", 21108 => "10011000", 21109 => "11111000", 21110 => "10110111", 21112 => "10000001", 21114 => "11011010", 21115 => "10110100", 21119 => "01000111", 21121 => "11110111", 21122 => "10100000", 21124 => "00110110", 21125 => "11111100", 21126 => "01011010", 21127 => "10001100", 21128 => "00100111", 21129 => "00111010", 21130 => "00111001", 21131 => "11011101", 21133 => "11110000", 21134 => "11111000", 21136 => "00000101", 21138 => "10111110", 21139 => "10110000", 21140 => "10101011", 21141 => "00100110", 21142 => "10101110", 21143 => "10011101", 21144 => "00110100", 21145 => "10010011", 21149 => "00011100", 21150 => "11000011", 21154 => "01001111", 21155 => "00001011", 21157 => "11010001", 21158 => "10110110", 21159 => "10000101", 21160 => "00010011", 21161 => "00110010", 21162 => "11111110", 21165 => "01001101", 21166 => "00111100", 21170 => "01000001", 21171 => "10001100", 21173 => "01101110", 21174 => "11111001", 21177 => "01101111", 21179 => "00110001", 21180 => "11011101", 21184 => "00100010", 21185 => "00001001", 21187 => "00110101", 21188 => "10100100", 21190 => "00000101", 21191 => "01110100", 21195 => "00111011", 21198 => "00111101", 21202 => "10110011", 21203 => "11010101", 21206 => "11111000", 21211 => "01110101", 21213 => "10111000", 21214 => "01111001", 21215 => "01011111", 21216 => "00001000", 21218 => "10010100", 21222 => "00111000", 21223 => "10111010", 21225 => "00111010", 21226 => "00110101", 21227 => "11011101", 21228 => "10111010", 21232 => "11111110", 21233 => "01101111", 21235 => "10111110", 21237 => "10110100", 21240 => "10111011", 21243 => "11110110", 21246 => "01010010", 21249 => "10000111", 21250 => "11000010", 21251 => "10011010", 21252 => "10010000", 21254 => "11000011", 21258 => "00101010", 21259 => "01100100", 21260 => "01111001", 21261 => "01110101", 21262 => "00010010", 21267 => "10110111", 21269 => "11001100", 21270 => "11101010", 21274 => "00000011", 21276 => "10000101", 21279 => "10001110", 21280 => "00111011", 21282 => "01100101", 21283 => "10001001", 21285 => "00100110", 21287 => "10100000", 21289 => "10000000", 21290 => "00001101", 21291 => "00010110", 21294 => "01111010", 21301 => "01111100", 21302 => "01101110", 21304 => "11111101", 21306 => "10010011", 21307 => "01100010", 21308 => "01100011", 21314 => "01101101", 21317 => "01110101", 21320 => "00011111", 21325 => "11001111", 21326 => "00111011", 21328 => "01010001", 21329 => "01110010", 21330 => "00110111", 21331 => "01100110", 21333 => "01101101", 21337 => "01110000", 21338 => "11100010", 21339 => "01010100", 21342 => "00001001", 21343 => "00011011", 21344 => "01100011", 21348 => "00100010", 21351 => "00110101", 21352 => "10011000", 21353 => "01110001", 21354 => "10111011", 21356 => "01110000", 21357 => "11111010", 21358 => "01100011", 21359 => "01111000", 21363 => "00111010", 21364 => "10111101", 21366 => "10011000", 21368 => "10000110", 21370 => "01011001", 21371 => "10010010", 21374 => "10100110", 21376 => "10000011", 21377 => "10100110", 21383 => "01011100", 21384 => "10010000", 21387 => "00101110", 21388 => "11000011", 21389 => "10111000", 21390 => "10001010", 21391 => "00110011", 21393 => "00100011", 21397 => "00010111", 21398 => "10111001", 21399 => "01010110", 21401 => "00010000", 21402 => "01111010", 21404 => "11100011", 21406 => "01011001", 21407 => "00111011", 21408 => "10111000", 21410 => "11110100", 21412 => "00001001", 21413 => "10110110", 21414 => "01000111", 21415 => "11001001", 21416 => "00100101", 21418 => "01101011", 21422 => "01010110", 21425 => "11110010", 21430 => "10010001", 21433 => "11100011", 21434 => "00000101", 21435 => "11100111", 21436 => "00011010", 21441 => "01010001", 21442 => "11000100", 21443 => "10011001", 21444 => "00000110", 21445 => "11011101", 21446 => "11100111", 21448 => "01011110", 21451 => "10000101", 21460 => "11100000", 21462 => "10000010", 21466 => "01001001", 21467 => "01111101", 21468 => "01000110", 21471 => "00111100", 21472 => "10110111", 21475 => "11110101", 21477 => "11101010", 21481 => "00111000", 21482 => "00111011", 21484 => "11110110", 21485 => "11111100", 21487 => "00011000", 21488 => "10001110", 21492 => "01111011", 21494 => "01010010", 21496 => "11101110", 21499 => "10010110", 21500 => "01010100", 21502 => "10101101", 21504 => "00100110", 21506 => "00010111", 21508 => "10001010", 21513 => "10000010", 21515 => "01000001", 21516 => "11100010", 21518 => "00111000", 21521 => "01011011", 21522 => "01011101", 21523 => "10111101", 21525 => "00001101", 21526 => "01101111", 21528 => "01100011", 21530 => "11111100", 21534 => "01110000", 21535 => "11011111", 21537 => "01101111", 21538 => "10001011", 21539 => "10111000", 21540 => "01011011", 21541 => "11001101", 21542 => "11000001", 21544 => "11100100", 21548 => "00111000", 21549 => "00100000", 21550 => "11101001", 21551 => "01110001", 21553 => "01000000", 21554 => "11001100", 21555 => "11101011", 21556 => "10011010", 21558 => "10011001", 21561 => "01110100", 21562 => "01011010", 21567 => "11110111", 21569 => "10101000", 21572 => "00011000", 21573 => "01001100", 21577 => "01110101", 21578 => "01000011", 21581 => "11011110", 21582 => "00110000", 21584 => "10010100", 21585 => "10011010", 21590 => "00000101", 21593 => "00110111", 21595 => "00010001", 21596 => "10100000", 21598 => "00111001", 21599 => "01010100", 21600 => "01011100", 21602 => "10110111", 21603 => "10011010", 21604 => "01110001", 21605 => "01000111", 21609 => "01101111", 21615 => "00001011", 21619 => "10100000", 21622 => "01000110", 21623 => "10001000", 21624 => "11100001", 21625 => "11101101", 21626 => "11110010", 21627 => "00100010", 21628 => "00100011", 21629 => "00111110", 21630 => "00101110", 21631 => "10011000", 21634 => "01011011", 21636 => "00000010", 21637 => "10110110", 21638 => "10011010", 21642 => "01100010", 21643 => "01111000", 21645 => "01101100", 21647 => "10011101", 21649 => "01111001", 21650 => "11111110", 21652 => "00110010", 21654 => "11001010", 21656 => "00110010", 21657 => "10100101", 21659 => "10111000", 21661 => "01001110", 21662 => "10101010", 21666 => "11111000", 21667 => "10010000", 21669 => "00011101", 21673 => "11111110", 21674 => "01101111", 21675 => "01010010", 21676 => "01010100", 21683 => "01000101", 21684 => "00100100", 21685 => "10010101", 21686 => "10110101", 21689 => "10110011", 21690 => "11111010", 21692 => "00100000", 21694 => "10010000", 21696 => "10010001", 21697 => "00101001", 21698 => "11011010", 21699 => "11000111", 21702 => "10000100", 21703 => "01101010", 21704 => "01100011", 21710 => "11001001", 21712 => "11011110", 21716 => "10111010", 21720 => "01010100", 21722 => "11111010", 21725 => "10001111", 21728 => "10000001", 21730 => "10110011", 21731 => "10101010", 21732 => "01101101", 21735 => "01010101", 21742 => "10100000", 21744 => "01010111", 21745 => "01001000", 21747 => "00000011", 21748 => "11110010", 21752 => "00010011", 21755 => "01110101", 21757 => "10000010", 21759 => "00111011", 21763 => "11001011", 21765 => "00001101", 21766 => "00000011", 21767 => "01100111", 21772 => "01001001", 21773 => "11001001", 21776 => "10010110", 21777 => "01000100", 21779 => "11110001", 21780 => "10111100", 21782 => "11011101", 21785 => "00100101", 21787 => "11100100", 21788 => "01001011", 21790 => "01101110", 21792 => "10111001", 21797 => "10001011", 21800 => "11111111", 21801 => "01100110", 21803 => "01010010", 21804 => "01010111", 21805 => "10001100", 21808 => "00110010", 21809 => "11010100", 21811 => "11100101", 21812 => "11111111", 21817 => "01011111", 21818 => "01111111", 21820 => "11100110", 21821 => "00010101", 21822 => "11011011", 21824 => "10110001", 21827 => "11111000", 21829 => "01111110", 21830 => "01011110", 21835 => "00001011", 21836 => "11110101", 21841 => "01111110", 21843 => "11111011", 21844 => "10100111", 21845 => "11000001", 21848 => "00110001", 21849 => "00010010", 21851 => "01010111", 21853 => "00101001", 21857 => "00010000", 21860 => "01100100", 21864 => "10101100", 21865 => "01001010", 21867 => "01010110", 21868 => "10100110", 21870 => "11010111", 21871 => "11101101", 21872 => "10110110", 21874 => "10100010", 21875 => "11111000", 21881 => "00011100", 21883 => "11101001", 21885 => "10001100", 21886 => "11010111", 21887 => "01010001", 21889 => "11111000", 21890 => "10111100", 21894 => "10000010", 21897 => "01111110", 21899 => "01110000", 21902 => "01100010", 21908 => "10111111", 21913 => "00101100", 21914 => "00110111", 21915 => "00101111", 21917 => "01001110", 21918 => "10101110", 21922 => "10000110", 21923 => "01111110", 21927 => "01001010", 21928 => "01101100", 21931 => "10001101", 21933 => "01111100", 21934 => "01011011", 21935 => "10010010", 21936 => "01000001", 21937 => "10010111", 21938 => "10100101", 21939 => "01000011", 21941 => "01111101", 21943 => "11110110", 21944 => "00100111", 21945 => "01011000", 21946 => "00101100", 21947 => "00000010", 21948 => "01100101", 21950 => "00000101", 21953 => "11001011", 21955 => "10000101", 21956 => "10101000", 21957 => "01010110", 21958 => "00110110", 21959 => "10010000", 21960 => "10101010", 21961 => "01000110", 21962 => "00101010", 21966 => "10111011", 21971 => "01010000", 21973 => "00111001", 21975 => "11101010", 21976 => "11011011", 21977 => "11111100", 21979 => "11110101", 21981 => "00010000", 21984 => "11110101", 21986 => "11101100", 21987 => "10000101", 21990 => "11010101", 21998 => "01001100", 22001 => "00111100", 22002 => "10100111", 22004 => "01111001", 22006 => "00101010", 22009 => "10110101", 22011 => "01100110", 22014 => "01100001", 22016 => "11110001", 22021 => "00101101", 22022 => "01110000", 22024 => "11100101", 22026 => "10110010", 22033 => "10001011", 22034 => "11000100", 22035 => "11110010", 22037 => "10010011", 22038 => "00101010", 22039 => "01001111", 22041 => "11000100", 22045 => "01011101", 22046 => "11110010", 22047 => "00100000", 22048 => "11000000", 22051 => "11110011", 22052 => "10101000", 22053 => "10110100", 22055 => "01010011", 22060 => "11011111", 22062 => "00100001", 22063 => "01001101", 22064 => "10111110", 22065 => "11000101", 22073 => "00001110", 22074 => "01101001", 22075 => "00100100", 22078 => "00100100", 22081 => "11100101", 22083 => "00001001", 22086 => "00010111", 22087 => "11000110", 22090 => "10110001", 22091 => "11100011", 22096 => "00111000", 22098 => "00100011", 22100 => "11111011", 22101 => "10111111", 22107 => "00110110", 22109 => "11111010", 22110 => "11001111", 22115 => "11111101", 22117 => "11101011", 22119 => "11010111", 22120 => "00101101", 22123 => "01111010", 22124 => "00100111", 22125 => "11011111", 22126 => "00010010", 22127 => "01010010", 22128 => "01100100", 22129 => "10111010", 22130 => "00100011", 22131 => "00100100", 22133 => "11010010", 22135 => "00011001", 22138 => "01101000", 22140 => "10010001", 22142 => "10000100", 22146 => "00100101", 22148 => "11111110", 22149 => "11111011", 22150 => "11110101", 22152 => "01011100", 22153 => "00001101", 22156 => "10100011", 22161 => "10101110", 22162 => "01011010", 22163 => "00100000", 22165 => "11111010", 22166 => "01100001", 22168 => "01111100", 22169 => "11100000", 22174 => "10010001", 22175 => "01001110", 22176 => "10101011", 22178 => "01011001", 22179 => "10101011", 22180 => "01101110", 22182 => "01011001", 22184 => "01000110", 22186 => "10111011", 22189 => "11011101", 22190 => "01110101", 22192 => "00111011", 22198 => "00001110", 22201 => "00111100", 22204 => "11010000", 22205 => "10111001", 22206 => "01011100", 22208 => "00100110", 22209 => "00001000", 22210 => "00001011", 22211 => "11000011", 22213 => "11111010", 22214 => "00000010", 22219 => "00111111", 22220 => "10001101", 22221 => "10000001", 22222 => "11001000", 22224 => "00100110", 22225 => "11001111", 22226 => "00100011", 22227 => "11010100", 22229 => "10100110", 22235 => "11001101", 22237 => "01111010", 22242 => "10111101", 22244 => "00110111", 22246 => "11001010", 22247 => "11110000", 22248 => "10110100", 22251 => "11011000", 22252 => "01100010", 22253 => "10111110", 22254 => "11010011", 22255 => "11011011", 22256 => "11101000", 22257 => "01001100", 22258 => "01101001", 22259 => "10101110", 22260 => "01101100", 22261 => "01001001", 22263 => "01101010", 22264 => "10010010", 22265 => "11101010", 22266 => "01110101", 22267 => "00000010", 22269 => "01110101", 22273 => "01100111", 22274 => "11110001", 22275 => "00100100", 22276 => "01011100", 22277 => "01110010", 22281 => "10110110", 22282 => "11000010", 22283 => "00100110", 22285 => "11010110", 22286 => "10110100", 22287 => "00100010", 22289 => "01011001", 22293 => "00111000", 22295 => "11110001", 22298 => "00000010", 22300 => "11010110", 22302 => "01010111", 22304 => "01000101", 22305 => "00001000", 22307 => "10111101", 22308 => "01110101", 22310 => "00000011", 22312 => "00001010", 22313 => "10110000", 22314 => "01110110", 22320 => "00010100", 22321 => "10111111", 22322 => "11111011", 22323 => "00111101", 22324 => "01110000", 22325 => "01100100", 22327 => "10110101", 22330 => "11000010", 22333 => "10001001", 22335 => "00001110", 22339 => "00010010", 22341 => "00001000", 22343 => "00111001", 22344 => "01001111", 22345 => "11000100", 22347 => "01111011", 22351 => "00000100", 22352 => "10000111", 22353 => "00000011", 22354 => "10011111", 22355 => "00000100", 22356 => "01111000", 22359 => "11100101", 22360 => "11010111", 22364 => "11011110", 22365 => "01100010", 22366 => "00010101", 22373 => "01100001", 22374 => "01010001", 22377 => "00110110", 22378 => "11000001", 22379 => "11000100", 22381 => "01111110", 22382 => "01100100", 22385 => "10111000", 22387 => "11111000", 22392 => "01011000", 22394 => "11101011", 22396 => "01110000", 22399 => "10010111", 22400 => "11111001", 22404 => "01101100", 22406 => "01010001", 22408 => "01010101", 22409 => "01000010", 22413 => "10101011", 22414 => "00101100", 22415 => "10101010", 22417 => "00110000", 22419 => "01110000", 22421 => "00000100", 22424 => "01111001", 22425 => "01111101", 22426 => "01010010", 22427 => "10000111", 22429 => "11111110", 22432 => "10110011", 22435 => "10101100", 22437 => "00010111", 22440 => "10010110", 22441 => "00011100", 22442 => "00111100", 22443 => "00010101", 22444 => "11001100", 22446 => "00001001", 22448 => "01111100", 22451 => "00110001", 22452 => "00110001", 22453 => "01110101", 22458 => "11000101", 22460 => "10110110", 22462 => "11011000", 22464 => "00011011", 22465 => "00011011", 22466 => "10010010", 22470 => "10101110", 22471 => "11011100", 22472 => "01110111", 22473 => "00111001", 22475 => "00100011", 22476 => "11110100", 22480 => "01001111", 22483 => "10001101", 22486 => "00010000", 22488 => "01110010", 22491 => "11100100", 22493 => "00001111", 22495 => "11110101", 22498 => "01001110", 22501 => "00011110", 22503 => "00000110", 22505 => "11000001", 22506 => "01111001", 22508 => "10111011", 22509 => "11000000", 22512 => "01111011", 22514 => "10100110", 22515 => "01011110", 22520 => "11100100", 22521 => "11011011", 22525 => "11101001", 22529 => "10010101", 22534 => "11001111", 22536 => "01100111", 22537 => "00001111", 22539 => "11111111", 22540 => "11111101", 22545 => "11101110", 22549 => "01010011", 22551 => "10010111", 22552 => "11011011", 22555 => "11110011", 22557 => "01000100", 22558 => "10110110", 22559 => "10011010", 22564 => "01000001", 22566 => "00111010", 22567 => "00100101", 22573 => "11000110", 22577 => "10001000", 22578 => "01111001", 22579 => "00010100", 22582 => "10001001", 22583 => "00010111", 22584 => "00111100", 22585 => "11111110", 22590 => "00010100", 22591 => "11001011", 22594 => "00000011", 22596 => "10111011", 22598 => "10110000", 22600 => "10101100", 22602 => "11000010", 22608 => "01011011", 22610 => "11001100", 22612 => "01100000", 22614 => "01101011", 22617 => "10001011", 22619 => "10010110", 22620 => "01111101", 22622 => "00011000", 22624 => "01110011", 22626 => "00110101", 22630 => "11011000", 22631 => "00100001", 22632 => "11011011", 22635 => "10000011", 22636 => "10111000", 22639 => "01101000", 22640 => "01011000", 22645 => "11111100", 22647 => "00100010", 22648 => "01101111", 22649 => "10010110", 22651 => "00100101", 22652 => "11001010", 22658 => "11101000", 22659 => "11011001", 22661 => "10110111", 22662 => "10100011", 22665 => "11111101", 22667 => "00100111", 22669 => "11000110", 22674 => "10000010", 22675 => "00001000", 22677 => "01111110", 22678 => "10110100", 22679 => "10101000", 22680 => "01110000", 22682 => "01101101", 22683 => "01100100", 22684 => "10000101", 22685 => "01100010", 22689 => "00000101", 22690 => "10110100", 22692 => "11000111", 22693 => "10111110", 22694 => "10101101", 22696 => "00010000", 22697 => "00101100", 22699 => "10000110", 22701 => "00001110", 22708 => "00100101", 22711 => "10000101", 22712 => "10100011", 22713 => "00110000", 22717 => "10011010", 22720 => "00001010", 22725 => "10001101", 22727 => "10110101", 22728 => "00001101", 22731 => "11010010", 22734 => "01011110", 22736 => "01011011", 22743 => "10000010", 22747 => "00011000", 22748 => "01011111", 22749 => "00011000", 22751 => "00101100", 22755 => "00111001", 22757 => "00110010", 22759 => "10001110", 22764 => "00011101", 22765 => "11011000", 22771 => "00111011", 22772 => "11110001", 22775 => "00100101", 22778 => "00100011", 22779 => "10111000", 22780 => "00001010", 22781 => "01011001", 22782 => "10000101", 22783 => "10011101", 22790 => "01110100", 22791 => "00111110", 22792 => "11010011", 22796 => "00110001", 22798 => "10101111", 22806 => "01101011", 22809 => "11101111", 22813 => "00010100", 22818 => "10010101", 22819 => "11000111", 22821 => "10110111", 22822 => "11101000", 22823 => "01000101", 22824 => "00000110", 22826 => "11011111", 22828 => "10011100", 22829 => "00011010", 22830 => "00010001", 22832 => "00011011", 22836 => "01001110", 22837 => "01111101", 22838 => "01100101", 22839 => "00001111", 22841 => "10001001", 22845 => "01000110", 22846 => "11010111", 22850 => "01100101", 22851 => "01101001", 22852 => "00001100", 22853 => "01011110", 22854 => "00011011", 22855 => "01011110", 22858 => "00100000", 22860 => "01010111", 22861 => "00010010", 22862 => "10111011", 22864 => "00011101", 22866 => "10011101", 22871 => "01100111", 22872 => "01101100", 22877 => "10100011", 22881 => "10101100", 22882 => "10110101", 22884 => "00001111", 22887 => "00111011", 22889 => "10010011", 22890 => "00111001", 22891 => "00000010", 22892 => "00011000", 22894 => "10010011", 22895 => "10111110", 22896 => "11011000", 22897 => "10010010", 22898 => "01111000", 22899 => "00111011", 22900 => "11000001", 22901 => "00010000", 22908 => "11100011", 22910 => "10011111", 22912 => "01001011", 22913 => "00110110", 22915 => "11001001", 22916 => "00010101", 22918 => "11101001", 22919 => "01011100", 22920 => "01100011", 22923 => "00011110", 22924 => "10111001", 22926 => "01001101", 22929 => "00111101", 22930 => "01110101", 22931 => "10100010", 22932 => "11110100", 22933 => "10111010", 22935 => "10111011", 22938 => "00110101", 22939 => "10100000", 22941 => "00000011", 22942 => "01111000", 22944 => "11001111", 22945 => "01100011", 22947 => "00101000", 22950 => "10111000", 22952 => "01101001", 22955 => "11100100", 22957 => "10110101", 22959 => "01100101", 22960 => "01111000", 22964 => "10101001", 22965 => "01110100", 22968 => "01010111", 22970 => "00000101", 22971 => "01100111", 22972 => "00011111", 22973 => "00001101", 22974 => "11000000", 22975 => "01100111", 22976 => "00110110", 22980 => "00110111", 22983 => "10000010", 22987 => "10100100", 22988 => "10001110", 22992 => "00101000", 22993 => "00110111", 22995 => "01000101", 22996 => "01100011", 22997 => "01101111", 22999 => "00111010", 23002 => "01001001", 23003 => "01100010", 23006 => "01000110", 23008 => "10101010", 23009 => "10001010", 23010 => "10000110", 23012 => "01110010", 23013 => "10111101", 23015 => "00101110", 23017 => "11110110", 23022 => "01110011", 23025 => "00110011", 23026 => "01011010", 23027 => "11101100", 23029 => "01100110", 23032 => "01001110", 23036 => "01010011", 23040 => "10001010", 23041 => "11011101", 23042 => "01000100", 23044 => "01101101", 23045 => "00010100", 23047 => "01101010", 23048 => "01000011", 23049 => "00100010", 23050 => "10010010", 23053 => "01101000", 23054 => "00011101", 23056 => "11000110", 23058 => "11101111", 23060 => "11111101", 23061 => "01111011", 23065 => "01111111", 23066 => "11111010", 23067 => "11000101", 23068 => "01001001", 23071 => "10101010", 23073 => "01110010", 23074 => "00101110", 23081 => "01100010", 23082 => "01101101", 23083 => "11001011", 23085 => "01111011", 23086 => "11100001", 23087 => "10001011", 23088 => "01100000", 23094 => "10000001", 23095 => "01110110", 23099 => "00101111", 23102 => "01000011", 23103 => "01011101", 23104 => "10001101", 23106 => "11001011", 23107 => "11110110", 23112 => "01111001", 23113 => "00001011", 23114 => "10001100", 23115 => "01001100", 23117 => "10011111", 23119 => "11001111", 23120 => "01000110", 23122 => "11110101", 23123 => "10001110", 23124 => "00000011", 23128 => "00111101", 23129 => "11110000", 23130 => "01011010", 23132 => "11000011", 23134 => "10011011", 23136 => "10000110", 23137 => "01110110", 23139 => "00011000", 23141 => "01111001", 23142 => "10110000", 23145 => "00101011", 23146 => "11000011", 23149 => "11100101", 23150 => "00100101", 23151 => "00010110", 23154 => "11001101", 23156 => "11100010", 23158 => "11111001", 23159 => "11010011", 23162 => "00101010", 23163 => "00010100", 23165 => "10110001", 23166 => "10110001", 23168 => "10001001", 23169 => "11110011", 23170 => "11111000", 23171 => "11011000", 23172 => "01001110", 23173 => "00000010", 23179 => "11100101", 23181 => "01001011", 23183 => "11001010", 23184 => "11011101", 23186 => "00001001", 23187 => "01010001", 23191 => "10001110", 23192 => "00100110", 23193 => "00001011", 23195 => "10110110", 23196 => "01110000", 23200 => "10011001", 23208 => "01101000", 23209 => "10100111", 23211 => "10000101", 23213 => "11000010", 23216 => "01011001", 23217 => "01111000", 23219 => "10001010", 23220 => "00010000", 23225 => "10101000", 23227 => "10101010", 23228 => "10010001", 23231 => "01100111", 23233 => "01000000", 23234 => "00111000", 23237 => "11011101", 23238 => "10111000", 23239 => "00111110", 23242 => "11001001", 23245 => "01000110", 23247 => "10111000", 23251 => "01010111", 23255 => "00111011", 23256 => "01110100", 23259 => "00110011", 23261 => "10010110", 23266 => "10010100", 23267 => "01101110", 23268 => "00110000", 23269 => "01100111", 23270 => "10011000", 23273 => "00101011", 23278 => "10101111", 23279 => "11111111", 23280 => "10011111", 23282 => "11000100", 23284 => "00101010", 23287 => "01101101", 23292 => "00000111", 23294 => "00100001", 23295 => "00111110", 23296 => "00100110", 23297 => "11111101", 23298 => "01011101", 23300 => "11000100", 23305 => "10011011", 23306 => "00001100", 23307 => "00011100", 23311 => "01001110", 23313 => "01011111", 23316 => "10111110", 23319 => "11010101", 23325 => "01101111", 23326 => "10110000", 23328 => "01011011", 23333 => "00011001", 23335 => "00110101", 23336 => "00100000", 23337 => "10001010", 23339 => "00011011", 23340 => "11001101", 23344 => "11001010", 23346 => "11000000", 23348 => "11000000", 23349 => "01011101", 23350 => "01000011", 23351 => "01011110", 23352 => "01001000", 23353 => "11100100", 23354 => "01110010", 23357 => "10100000", 23359 => "01011100", 23368 => "01001111", 23369 => "00100100", 23370 => "11101000", 23371 => "00000110", 23372 => "01100110", 23373 => "10000111", 23376 => "11100000", 23380 => "01011111", 23381 => "01011100", 23382 => "11010010", 23383 => "01000111", 23384 => "11111010", 23387 => "10101111", 23392 => "01010000", 23394 => "01001001", 23395 => "10000010", 23396 => "01000001", 23397 => "10011001", 23398 => "01011100", 23399 => "11110011", 23402 => "11010101", 23407 => "11100100", 23408 => "11110100", 23409 => "01100000", 23413 => "10011101", 23414 => "10100011", 23416 => "10000011", 23417 => "00010111", 23418 => "00101010", 23419 => "10111111", 23420 => "01011100", 23422 => "10010101", 23423 => "11001101", 23424 => "11100100", 23425 => "10011100", 23426 => "00010001", 23429 => "10101100", 23430 => "01101110", 23431 => "01101100", 23432 => "00110100", 23434 => "00101110", 23435 => "01011100", 23437 => "10001011", 23439 => "01010111", 23442 => "01101101", 23445 => "10010101", 23446 => "01001100", 23447 => "10010010", 23449 => "01101010", 23450 => "10011000", 23451 => "00011111", 23452 => "01100111", 23453 => "10100011", 23455 => "10101000", 23456 => "11000011", 23459 => "11010010", 23461 => "00101111", 23467 => "01010111", 23469 => "00011101", 23474 => "10111000", 23478 => "00011010", 23479 => "10101010", 23480 => "10101001", 23481 => "01110000", 23484 => "01111000", 23486 => "00101001", 23487 => "00110000", 23490 => "10010011", 23492 => "10001101", 23493 => "10001100", 23495 => "11110100", 23496 => "01011011", 23502 => "10010010", 23504 => "10100000", 23510 => "11100101", 23511 => "10001010", 23512 => "10111110", 23514 => "01111100", 23516 => "10011111", 23518 => "10100000", 23519 => "10101110", 23521 => "10110011", 23523 => "00111011", 23524 => "10010101", 23525 => "11000110", 23526 => "11101111", 23528 => "11000111", 23531 => "11110101", 23535 => "10101100", 23536 => "10011101", 23537 => "01001111", 23538 => "00011000", 23539 => "00011111", 23540 => "01001000", 23541 => "11111010", 23543 => "10100001", 23544 => "11001011", 23546 => "11000111", 23548 => "11100100", 23549 => "11101111", 23552 => "11110001", 23555 => "00010111", 23558 => "00000110", 23563 => "01111010", 23565 => "11111101", 23567 => "01110110", 23568 => "00010110", 23569 => "11011110", 23573 => "11100011", 23576 => "01110001", 23577 => "01100110", 23579 => "00110001", 23581 => "10011010", 23582 => "11010001", 23588 => "10011101", 23589 => "10100001", 23590 => "00000001", 23596 => "01110001", 23598 => "11000101", 23599 => "00101111", 23604 => "10100010", 23606 => "01100111", 23607 => "10011011", 23616 => "01010111", 23618 => "00101001", 23619 => "01111101", 23620 => "11100100", 23621 => "00001101", 23623 => "01001010", 23624 => "00010101", 23627 => "01000010", 23629 => "10000100", 23632 => "00101110", 23633 => "11110000", 23638 => "01001100", 23639 => "00101100", 23640 => "00101101", 23642 => "01000101", 23643 => "11110000", 23645 => "10000100", 23646 => "00110000", 23647 => "10010111", 23650 => "10001011", 23651 => "11000011", 23652 => "01101111", 23653 => "00110011", 23655 => "10001100", 23656 => "10001011", 23657 => "01101010", 23658 => "01000111", 23659 => "10100101", 23660 => "01110110", 23661 => "01001101", 23662 => "10110011", 23668 => "00101100", 23670 => "00001100", 23673 => "01000000", 23674 => "10011001", 23675 => "10010110", 23677 => "00011000", 23678 => "11110110", 23679 => "01101101", 23680 => "11010101", 23683 => "10001100", 23684 => "00000011", 23686 => "11101111", 23687 => "11011011", 23691 => "11011100", 23692 => "10110010", 23693 => "01110110", 23697 => "10111010", 23699 => "00001011", 23700 => "01100011", 23701 => "10111111", 23703 => "11000111", 23707 => "01111000", 23713 => "01000101", 23714 => "11101111", 23719 => "01001111", 23720 => "01100110", 23721 => "11101011", 23726 => "00101010", 23730 => "01110011", 23731 => "01101101", 23732 => "00011011", 23733 => "10010100", 23736 => "11110111", 23738 => "01000011", 23739 => "01011011", 23741 => "01101000", 23743 => "11100111", 23745 => "11000101", 23747 => "01011001", 23749 => "11001101", 23751 => "10000010", 23755 => "10001010", 23759 => "11001010", 23760 => "10011100", 23761 => "11011010", 23763 => "00010000", 23773 => "00111111", 23775 => "01110101", 23776 => "10010011", 23777 => "10100111", 23778 => "00101100", 23779 => "01101100", 23780 => "10100001", 23781 => "00111011", 23785 => "01000110", 23786 => "11101100", 23787 => "01001101", 23792 => "01100111", 23795 => "00001010", 23798 => "01100010", 23799 => "10010000", 23800 => "11000111", 23802 => "00010100", 23809 => "10110001", 23812 => "00011111", 23813 => "01010101", 23816 => "11011001", 23817 => "10111000", 23821 => "10100000", 23822 => "00100010", 23823 => "11000011", 23824 => "11000111", 23825 => "00101110", 23828 => "00101011", 23829 => "00100010", 23830 => "00110100", 23831 => "10000000", 23832 => "10111010", 23834 => "01010110", 23838 => "11110011", 23839 => "00010111", 23842 => "01010100", 23843 => "00000010", 23847 => "10001100", 23848 => "01100001", 23851 => "10010001", 23854 => "00101100", 23857 => "00100111", 23859 => "00000010", 23860 => "11110011", 23861 => "10010010", 23864 => "00110100", 23865 => "11100010", 23866 => "10000010", 23867 => "00010001", 23868 => "01000110", 23869 => "10111111", 23870 => "01010110", 23874 => "01100111", 23875 => "01011001", 23876 => "00111001", 23877 => "11100101", 23880 => "10010100", 23881 => "10000111", 23882 => "11110111", 23886 => "11000000", 23887 => "10001101", 23888 => "01100000", 23891 => "01011101", 23893 => "00100101", 23894 => "10001110", 23897 => "00110101", 23899 => "11101111", 23902 => "00101011", 23904 => "00110100", 23905 => "01000001", 23908 => "11100110", 23910 => "00011000", 23911 => "00001000", 23913 => "10100101", 23914 => "11111000", 23915 => "00001111", 23916 => "00101100", 23923 => "10101110", 23924 => "01011111", 23926 => "10111000", 23930 => "00001000", 23935 => "10110011", 23937 => "11110111", 23938 => "01011011", 23939 => "11100001", 23940 => "00011100", 23942 => "10110100", 23943 => "00101001", 23946 => "11011000", 23947 => "11000110", 23950 => "10010110", 23952 => "11010111", 23954 => "11011110", 23957 => "10011001", 23961 => "01010101", 23963 => "10111100", 23964 => "01100110", 23965 => "00110001", 23969 => "01111011", 23970 => "01001111", 23971 => "10000110", 23972 => "00100100", 23974 => "01101101", 23975 => "00111011", 23977 => "10001100", 23978 => "10001000", 23980 => "00110100", 23981 => "10111111", 23983 => "11011011", 23984 => "00111001", 23985 => "11100001", 23986 => "01100000", 23988 => "11001100", 23990 => "10100100", 23991 => "10110110", 23992 => "10111011", 23993 => "00100100", 23995 => "10001011", 23997 => "11000010", 24001 => "10000111", 24002 => "01101010", 24003 => "01101100", 24004 => "11001011", 24005 => "01010011", 24007 => "01100111", 24008 => "01110000", 24011 => "00001111", 24021 => "10000010", 24023 => "11101100", 24025 => "00010011", 24027 => "01100000", 24028 => "01100111", 24030 => "10011110", 24031 => "10001101", 24033 => "10100101", 24034 => "11101011", 24036 => "01011001", 24039 => "10000100", 24042 => "11101011", 24043 => "01011011", 24047 => "01100101", 24054 => "01001101", 24059 => "11110010", 24060 => "11011101", 24061 => "00100110", 24062 => "00101101", 24063 => "11110110", 24064 => "00111001", 24069 => "11111111", 24070 => "10001000", 24071 => "10110101", 24072 => "00011000", 24073 => "00110101", 24075 => "10110100", 24076 => "11100100", 24078 => "01000000", 24080 => "00101100", 24081 => "01011000", 24082 => "10111001", 24085 => "10011000", 24086 => "00111011", 24089 => "10101011", 24090 => "11000101", 24092 => "10100011", 24096 => "01001100", 24099 => "11000001", 24100 => "11110100", 24101 => "00011110", 24102 => "10010010", 24105 => "01100010", 24109 => "11000011", 24113 => "11000011", 24117 => "10001101", 24118 => "01001000", 24121 => "10000111", 24124 => "00111011", 24126 => "00111100", 24127 => "00001110", 24128 => "01100011", 24132 => "01111011", 24134 => "00010101", 24136 => "01100011", 24137 => "00010111", 24139 => "00110100", 24140 => "11000001", 24141 => "00111100", 24142 => "00011001", 24143 => "10101110", 24146 => "00110000", 24148 => "10011000", 24149 => "10101100", 24150 => "11100111", 24158 => "00110001", 24159 => "11101011", 24161 => "10011010", 24162 => "10001000", 24163 => "10010110", 24165 => "11000000", 24171 => "01000010", 24173 => "11000011", 24175 => "01101111", 24176 => "01100001", 24177 => "00101100", 24178 => "11101110", 24180 => "10001011", 24184 => "10111110", 24186 => "11000101", 24189 => "00100000", 24191 => "10101101", 24192 => "10011011", 24194 => "01010111", 24195 => "00101000", 24197 => "00101101", 24198 => "00010010", 24199 => "01111010", 24200 => "00101100", 24204 => "01001010", 24205 => "10000001", 24207 => "11010001", 24210 => "00111110", 24212 => "11001000", 24214 => "01111111", 24215 => "01010011", 24216 => "00111001", 24217 => "00110000", 24218 => "10000001", 24222 => "00000010", 24224 => "10110111", 24225 => "11011110", 24230 => "01000001", 24237 => "00010100", 24240 => "01100011", 24245 => "00010100", 24246 => "00110011", 24248 => "11011001", 24249 => "00010100", 24252 => "11101010", 24254 => "01100000", 24255 => "00011101", 24259 => "00000100", 24263 => "00000010", 24266 => "10010000", 24270 => "10010011", 24271 => "11000111", 24272 => "01011001", 24275 => "10001100", 24276 => "10001001", 24279 => "11101101", 24282 => "11000000", 24284 => "00110001", 24285 => "00011000", 24286 => "11001101", 24287 => "01001010", 24288 => "11111001", 24291 => "00010110", 24293 => "11101001", 24295 => "00010101", 24296 => "11001011", 24298 => "11100100", 24301 => "11011000", 24302 => "00010000", 24305 => "01101001", 24307 => "11110000", 24308 => "01011000", 24309 => "10001101", 24315 => "11011101", 24320 => "11110011", 24321 => "11111010", 24323 => "01001100", 24325 => "10100111", 24326 => "01110111", 24329 => "10101010", 24330 => "11100111", 24331 => "00101010", 24333 => "00010101", 24334 => "00000001", 24336 => "00101111", 24337 => "01011000", 24338 => "11100101", 24341 => "01100000", 24342 => "00001000", 24344 => "11001110", 24345 => "11000101", 24346 => "11111100", 24347 => "01110011", 24348 => "01101000", 24349 => "00100111", 24350 => "11001101", 24356 => "10011000", 24357 => "11111100", 24359 => "10011100", 24360 => "11110000", 24361 => "00100011", 24362 => "11010010", 24365 => "00011100", 24367 => "10110111", 24368 => "11010010", 24369 => "00011111", 24371 => "00111101", 24374 => "01100111", 24375 => "01001000", 24377 => "01000000", 24378 => "00100111", 24381 => "10111110", 24382 => "00001111", 24383 => "11110011", 24384 => "10011110", 24385 => "01010001", 24386 => "11110011", 24389 => "10110000", 24391 => "11001110", 24393 => "00110001", 24395 => "00110100", 24396 => "11001110", 24398 => "00001010", 24399 => "11101100", 24401 => "10101101", 24402 => "10001110", 24403 => "00000111", 24406 => "01011111", 24407 => "10110011", 24408 => "01011000", 24409 => "00110000", 24414 => "01100001", 24415 => "11100111", 24416 => "00000001", 24417 => "11010111", 24422 => "10101110", 24426 => "11110000", 24429 => "01110011", 24431 => "10000101", 24438 => "00001100", 24440 => "01001011", 24441 => "11001001", 24442 => "00100001", 24443 => "10111001", 24444 => "00110010", 24446 => "01001110", 24447 => "00110101", 24448 => "11011100", 24449 => "01110010", 24450 => "00001011", 24451 => "01011001", 24452 => "01000000", 24453 => "10000000", 24454 => "01110001", 24455 => "01000100", 24456 => "11000001", 24457 => "10001110", 24459 => "10011111", 24463 => "10100010", 24465 => "10010101", 24466 => "11010000", 24467 => "00001111", 24469 => "00111101", 24470 => "00001000", 24472 => "11100101", 24474 => "00010010", 24475 => "01001111", 24476 => "11011011", 24478 => "00010001", 24479 => "01101100", 24480 => "01010000", 24481 => "11100110", 24482 => "01010010", 24483 => "01010010", 24484 => "01110000", 24487 => "01001101", 24488 => "01001010", 24490 => "11010101", 24491 => "00011001", 24495 => "00010011", 24499 => "11001011", 24500 => "11101010", 24501 => "11001101", 24502 => "01000111", 24503 => "11010001", 24506 => "10000110", 24509 => "10000110", 24510 => "00001110", 24511 => "11000110", 24515 => "10110010", 24519 => "00111101", 24521 => "11101101", 24523 => "11000111", 24524 => "00100100", 24526 => "10110101", 24527 => "01000000", 24531 => "10001010", 24532 => "10110111", 24534 => "11101101", 24535 => "11110001", 24536 => "10111001", 24538 => "10111101", 24542 => "11000111", 24543 => "10100110", 24546 => "11000101", 24548 => "00101100", 24549 => "11101100", 24551 => "00101111", 24553 => "00110001", 24554 => "00110000", 24558 => "11111111", 24560 => "11110000", 24561 => "01111010", 24563 => "10011010", 24565 => "01011101", 24567 => "10011111", 24568 => "00110000", 24572 => "01100110", 24573 => "01111001", 24576 => "10110010", 24577 => "11100101", 24578 => "00000001", 24580 => "00101100", 24583 => "01010101", 24584 => "11110101", 24585 => "11011011", 24587 => "00110001", 24592 => "00100001", 24593 => "01000110", 24594 => "11000111", 24597 => "01000000", 24598 => "11011111", 24599 => "11100000", 24600 => "10000110", 24602 => "11000001", 24603 => "10111110", 24604 => "01001000", 24605 => "10011001", 24610 => "00100110", 24611 => "01000001", 24612 => "01001011", 24613 => "10010100", 24616 => "11110110", 24618 => "11111110", 24623 => "00010010", 24624 => "11100001", 24627 => "00010110", 24629 => "10101000", 24631 => "00011100", 24634 => "11010011", 24635 => "11010011", 24637 => "11111100", 24639 => "10001010", 24646 => "10111101", 24649 => "01000010", 24651 => "01001111", 24652 => "11100110", 24653 => "11100010", 24655 => "00011111", 24656 => "11000011", 24661 => "01001001", 24664 => "10110110", 24665 => "00011001", 24670 => "11000100", 24672 => "10100100", 24675 => "01011000", 24678 => "00010001", 24680 => "11000111", 24685 => "10101001", 24687 => "10001111", 24689 => "11010011", 24690 => "01011110", 24693 => "10001000", 24694 => "10101011", 24695 => "10000011", 24697 => "00001111", 24700 => "01100011", 24701 => "10100011", 24706 => "01111000", 24707 => "00011011", 24708 => "00001111", 24709 => "00100010", 24710 => "00001000", 24711 => "10001111", 24715 => "01110111", 24716 => "00101000", 24717 => "00100110", 24719 => "10000101", 24722 => "00101110", 24723 => "11010000", 24724 => "01001110", 24725 => "01111100", 24727 => "11010001", 24728 => "10000010", 24729 => "00110111", 24731 => "10111111", 24733 => "00011101", 24734 => "00011011", 24735 => "11000100", 24737 => "11100001", 24738 => "10010111", 24740 => "00001101", 24741 => "00000100", 24742 => "10101000", 24745 => "01100100", 24746 => "10111001", 24748 => "00001010", 24749 => "11001011", 24750 => "11001011", 24751 => "10101101", 24754 => "00010001", 24755 => "01101100", 24756 => "11100100", 24759 => "01010010", 24761 => "11010101", 24763 => "10111010", 24766 => "00100010", 24770 => "00000101", 24771 => "01001011", 24775 => "10100001", 24777 => "11100101", 24779 => "01111011", 24781 => "11110101", 24782 => "01000110", 24784 => "10011010", 24789 => "11100101", 24790 => "01110010", 24791 => "00010101", 24792 => "10000100", 24794 => "00110100", 24796 => "11000010", 24797 => "00010001", 24798 => "10001011", 24800 => "10111100", 24801 => "10101010", 24802 => "10110000", 24808 => "01101011", 24809 => "00010110", 24810 => "00001110", 24811 => "11101000", 24816 => "11001100", 24817 => "11000111", 24819 => "01111011", 24820 => "10110111", 24821 => "01000000", 24823 => "10110110", 24825 => "10010000", 24829 => "01001000", 24830 => "00111000", 24831 => "01101011", 24833 => "10011000", 24835 => "00101100", 24837 => "10011100", 24838 => "01011101", 24842 => "01110001", 24844 => "01010010", 24846 => "11010100", 24848 => "11000110", 24849 => "11110000", 24854 => "10101000", 24857 => "11011110", 24861 => "11110011", 24862 => "11101010", 24864 => "01001111", 24867 => "00111100", 24873 => "11110001", 24874 => "11011011", 24876 => "10001000", 24877 => "11101111", 24878 => "01111111", 24879 => "01101010", 24882 => "10000100", 24887 => "00001110", 24888 => "11110010", 24889 => "11000000", 24890 => "00010001", 24894 => "10100110", 24897 => "11001001", 24900 => "00000111", 24901 => "10001001", 24902 => "11111110", 24905 => "11011011", 24906 => "00110101", 24907 => "01001101", 24908 => "01100011", 24913 => "01101101", 24915 => "01001010", 24916 => "11010000", 24917 => "10100010", 24918 => "11011000", 24919 => "00011101", 24926 => "00111011", 24931 => "00110101", 24932 => "00010000", 24933 => "00111011", 24934 => "00110111", 24935 => "01110111", 24939 => "01101010", 24942 => "01111110", 24943 => "01010010", 24945 => "00100101", 24948 => "10100001", 24950 => "01100001", 24951 => "01100110", 24952 => "01100001", 24953 => "11110100", 24955 => "00001110", 24961 => "11010111", 24962 => "01101100", 24963 => "10111100", 24964 => "10101000", 24965 => "00111110", 24972 => "00101110", 24976 => "00111011", 24978 => "10011010", 24979 => "11100111", 24980 => "01011001", 24985 => "10000101", 24986 => "01001001", 24988 => "11010110", 24989 => "11100110", 24993 => "11111110", 24995 => "00011101", 24999 => "11010011", 25000 => "10001100", 25002 => "00001010", 25005 => "11100000", 25006 => "11001111", 25007 => "00111001", 25008 => "01010001", 25012 => "01011001", 25015 => "01110110", 25017 => "00111000", 25019 => "11110000", 25022 => "01110001", 25023 => "01111101", 25025 => "01111101", 25029 => "11101011", 25031 => "00100101", 25034 => "10111101", 25036 => "11100001", 25037 => "00101001", 25039 => "10001010", 25042 => "00011010", 25043 => "01110111", 25045 => "10000010", 25047 => "01001101", 25048 => "11011100", 25050 => "11111110", 25051 => "01010111", 25052 => "01101001", 25054 => "01101110", 25058 => "00100011", 25060 => "00000111", 25061 => "00111110", 25062 => "11011011", 25064 => "00011011", 25067 => "11101000", 25068 => "10010100", 25069 => "01000111", 25070 => "10110001", 25072 => "01111111", 25074 => "11010010", 25075 => "10100011", 25082 => "00001100", 25083 => "01110010", 25088 => "01100000", 25089 => "10100110", 25091 => "10100100", 25093 => "01010111", 25095 => "10000011", 25097 => "01101011", 25098 => "11101000", 25100 => "11010001", 25101 => "10111110", 25104 => "01110110", 25106 => "10100010", 25109 => "10000001", 25110 => "00111101", 25111 => "10010100", 25113 => "01001101", 25114 => "11101100", 25116 => "01000111", 25121 => "10110110", 25123 => "11010000", 25125 => "00101000", 25128 => "00101000", 25129 => "01111000", 25132 => "10000011", 25133 => "01111000", 25135 => "00101001", 25136 => "10010101", 25138 => "10001111", 25140 => "11001010", 25142 => "00001010", 25143 => "00000011", 25144 => "00011010", 25145 => "00001101", 25148 => "01011000", 25149 => "01111000", 25150 => "01010101", 25153 => "00110000", 25155 => "11011101", 25156 => "11100001", 25159 => "10000001", 25161 => "11010000", 25162 => "11101010", 25163 => "00101000", 25167 => "00110110", 25169 => "11001001", 25175 => "00111110", 25176 => "01110010", 25177 => "00011110", 25179 => "01011001", 25181 => "11100111", 25182 => "10010111", 25183 => "00110111", 25184 => "01001010", 25185 => "01100100", 25187 => "11100101", 25188 => "10001110", 25190 => "00111001", 25191 => "00110101", 25192 => "10101101", 25193 => "10100000", 25194 => "10011100", 25199 => "00000111", 25201 => "11111111", 25205 => "11010100", 25207 => "01010100", 25208 => "11010110", 25210 => "00111000", 25212 => "11001101", 25214 => "01001110", 25215 => "00110011", 25216 => "01001111", 25217 => "01110000", 25219 => "01100011", 25221 => "10100111", 25222 => "01011010", 25225 => "11001110", 25231 => "01111011", 25232 => "00111110", 25233 => "11000110", 25234 => "00000010", 25237 => "01101110", 25239 => "00001110", 25240 => "10000110", 25241 => "11000001", 25242 => "00100001", 25243 => "10000001", 25245 => "00111010", 25248 => "00010010", 25249 => "11001011", 25250 => "01110011", 25251 => "01111011", 25252 => "11011010", 25254 => "10001100", 25257 => "11111010", 25258 => "00110111", 25261 => "00000110", 25269 => "11110111", 25271 => "00001000", 25272 => "11010000", 25273 => "10111001", 25274 => "00001100", 25275 => "01010011", 25276 => "11000110", 25279 => "11100011", 25281 => "10000100", 25282 => "00110001", 25283 => "00101100", 25289 => "11001110", 25292 => "10110011", 25293 => "10010100", 25294 => "00001110", 25295 => "01001110", 25296 => "00110010", 25297 => "10011110", 25302 => "10001101", 25303 => "01100101", 25306 => "00110111", 25309 => "11100010", 25310 => "01011010", 25313 => "11111100", 25314 => "01111001", 25315 => "10101011", 25316 => "00101000", 25319 => "00010111", 25320 => "10001001", 25321 => "10000010", 25322 => "00100001", 25323 => "01110100", 25327 => "10100000", 25330 => "01101101", 25334 => "11100111", 25337 => "01110001", 25338 => "11011011", 25340 => "11010000", 25341 => "00100011", 25342 => "11110010", 25346 => "00001010", 25347 => "01000101", 25348 => "00001100", 25349 => "00110101", 25352 => "01010111", 25356 => "01111111", 25357 => "01111111", 25358 => "10100000", 25359 => "11011100", 25361 => "01010100", 25364 => "00101100", 25365 => "10100100", 25369 => "10000011", 25370 => "01111101", 25371 => "01011110", 25375 => "10110110", 25378 => "11000100", 25382 => "11101011", 25383 => "01100011", 25385 => "10111010", 25386 => "00001001", 25388 => "11110010", 25390 => "10010000", 25391 => "11010101", 25392 => "01000000", 25395 => "11100001", 25398 => "11010100", 25403 => "11110011", 25406 => "11110100", 25409 => "01101001", 25410 => "00011010", 25411 => "01001000", 25413 => "10100011", 25414 => "01000111", 25415 => "01011000", 25417 => "00001111", 25419 => "11001110", 25420 => "00101010", 25421 => "01101010", 25424 => "11110000", 25425 => "10000000", 25426 => "01111010", 25428 => "11100011", 25429 => "10101001", 25433 => "10110001", 25434 => "01000110", 25438 => "00001100", 25440 => "00101011", 25442 => "10000100", 25443 => "01100111", 25444 => "00010001", 25449 => "11011111", 25450 => "10101000", 25451 => "11110101", 25452 => "01000011", 25455 => "00100101", 25458 => "10111000", 25459 => "10010101", 25460 => "10001100", 25464 => "10010100", 25465 => "11001111", 25466 => "11110110", 25469 => "00000010", 25470 => "11001110", 25471 => "11000011", 25474 => "10001001", 25481 => "00011110", 25487 => "11101000", 25488 => "01111110", 25489 => "11100110", 25490 => "01011011", 25491 => "10011101", 25493 => "00001111", 25494 => "11111000", 25495 => "11100100", 25497 => "01010110", 25498 => "11110010", 25503 => "01011011", 25504 => "11000010", 25506 => "00101011", 25507 => "11011110", 25509 => "00100101", 25513 => "11111000", 25515 => "11000011", 25520 => "10001111", 25523 => "01001111", 25524 => "00111110", 25525 => "11110011", 25527 => "01001001", 25528 => "00100100", 25530 => "10000001", 25534 => "00101011", 25535 => "10101000", 25538 => "11000000", 25539 => "10010110", 25540 => "11111000", 25546 => "01010111", 25547 => "10111111", 25550 => "11001100", 25551 => "01001100", 25554 => "00001110", 25555 => "11011111", 25556 => "10011100", 25559 => "10011000", 25560 => "01111011", 25562 => "01110010", 25563 => "10111100", 25565 => "00000110", 25567 => "11111011", 25569 => "11101101", 25570 => "00001101", 25573 => "01011000", 25578 => "10000100", 25580 => "10101000", 25582 => "00100101", 25584 => "11010011", 25585 => "00100111", 25588 => "01000001", 25590 => "10011110", 25591 => "01001010", 25593 => "01010011", 25594 => "01100001", 25596 => "00011001", 25598 => "10100011", 25599 => "00111011", 25600 => "11101110", 25601 => "11011010", 25603 => "01001110", 25604 => "10010000", 25605 => "11010001", 25607 => "00100011", 25608 => "01101000", 25609 => "10001001", 25610 => "01001111", 25611 => "11100111", 25612 => "00111011", 25613 => "11101110", 25614 => "11000111", 25615 => "01111011", 25616 => "11001000", 25618 => "10101010", 25620 => "11101110", 25621 => "10100000", 25622 => "10101101", 25625 => "10000011", 25626 => "00011000", 25627 => "10010000", 25628 => "00000110", 25629 => "11101110", 25630 => "00100011", 25631 => "01111011", 25633 => "00110111", 25635 => "00000110", 25636 => "01001100", 25639 => "00001100", 25642 => "01011001", 25643 => "00010010", 25648 => "11011110", 25653 => "00011100", 25655 => "11110000", 25656 => "01010011", 25659 => "01010000", 25660 => "11100011", 25662 => "10011010", 25663 => "11110100", 25667 => "01000011", 25672 => "00100000", 25676 => "11010100", 25679 => "10000110", 25682 => "10111101", 25684 => "11111000", 25686 => "01001110", 25687 => "11100000", 25689 => "11101111", 25690 => "10100100", 25692 => "10000111", 25693 => "00111111", 25694 => "10110100", 25695 => "10110011", 25698 => "01100011", 25700 => "10100011", 25701 => "01000100", 25702 => "10111011", 25704 => "00100011", 25706 => "00000001", 25707 => "00011011", 25709 => "00100010", 25713 => "01101110", 25718 => "10101101", 25719 => "00011000", 25721 => "01100011", 25723 => "10111000", 25724 => "10101001", 25725 => "11001101", 25726 => "01111000", 25728 => "10111011", 25729 => "10000110", 25730 => "00110110", 25732 => "01110010", 25733 => "10101110", 25734 => "11101101", 25736 => "11000100", 25737 => "01111111", 25740 => "00010111", 25742 => "01110100", 25743 => "01010000", 25746 => "01011111", 25751 => "01000101", 25755 => "01101110", 25756 => "11010101", 25758 => "01010010", 25760 => "10010100", 25761 => "01101111", 25763 => "00100000", 25764 => "10010110", 25766 => "00001010", 25768 => "11100111", 25770 => "01110011", 25772 => "11111010", 25773 => "01010010", 25774 => "01011111", 25775 => "01000100", 25778 => "10111111", 25779 => "00110110", 25782 => "01111000", 25783 => "00100001", 25784 => "10010100", 25787 => "00111111", 25788 => "10011010", 25789 => "00000101", 25790 => "00101010", 25791 => "01100110", 25793 => "01111011", 25794 => "00011000", 25797 => "11011001", 25799 => "01111000", 25806 => "01101110", 25807 => "10010111", 25808 => "11011000", 25809 => "10001111", 25810 => "10010010", 25811 => "11111001", 25812 => "00110111", 25816 => "01110101", 25818 => "10101011", 25820 => "01111110", 25823 => "10000011", 25825 => "11010011", 25826 => "01111000", 25827 => "00010011", 25830 => "01011011", 25833 => "11010000", 25835 => "00000101", 25836 => "01011100", 25838 => "10100110", 25839 => "10110001", 25841 => "10100111", 25843 => "10110110", 25849 => "00101000", 25850 => "10001110", 25851 => "10100001", 25852 => "10111010", 25854 => "01110011", 25855 => "11010100", 25862 => "00100111", 25863 => "00010000", 25864 => "10111100", 25867 => "10010011", 25869 => "11101011", 25870 => "01000010", 25873 => "11100011", 25875 => "11111111", 25876 => "01010100", 25877 => "00100010", 25879 => "01101100", 25883 => "01101100", 25887 => "11110011", 25890 => "10011100", 25892 => "00011110", 25893 => "10101001", 25898 => "00001011", 25899 => "10101000", 25900 => "00010010", 25901 => "01111100", 25903 => "11000110", 25904 => "01000110", 25910 => "00011000", 25911 => "00110100", 25912 => "00101010", 25913 => "00011001", 25914 => "00111000", 25917 => "01010000", 25919 => "10001101", 25920 => "11001011", 25921 => "01100101", 25923 => "01000000", 25924 => "00100011", 25926 => "01010101", 25928 => "01011011", 25931 => "00101110", 25937 => "10001101", 25939 => "00110010", 25943 => "00110111", 25946 => "10101001", 25948 => "01111101", 25949 => "10011010", 25950 => "00100111", 25951 => "00011111", 25952 => "00011011", 25953 => "00101001", 25954 => "10001100", 25955 => "10111001", 25957 => "11100101", 25959 => "10011100", 25960 => "01001010", 25962 => "00110100", 25964 => "11011000", 25966 => "11110100", 25968 => "10111000", 25969 => "01011010", 25973 => "01101010", 25976 => "11110101", 25977 => "00110101", 25979 => "10000101", 25980 => "01100100", 25982 => "00000101", 25986 => "11011111", 25988 => "01100100", 25989 => "01001111", 25991 => "10101110", 25993 => "00000001", 25995 => "11111000", 25996 => "01000101", 25997 => "00110100", 25998 => "01010110", 25999 => "00001101", 26001 => "10111101", 26004 => "00111101", 26007 => "10000110", 26008 => "01111011", 26009 => "11001001", 26010 => "10111010", 26012 => "11101110", 26013 => "11101111", 26014 => "00110000", 26017 => "11101000", 26018 => "00101101", 26019 => "00111010", 26021 => "00100100", 26024 => "10110111", 26028 => "01101011", 26029 => "11000110", 26032 => "10111010", 26034 => "10010101", 26038 => "11100010", 26039 => "00101111", 26044 => "10101100", 26046 => "00110101", 26047 => "11100101", 26049 => "01111110", 26051 => "00010010", 26056 => "01001000", 26059 => "01101000", 26062 => "10011010", 26063 => "01101011", 26064 => "10101110", 26065 => "01001000", 26069 => "11011001", 26070 => "01010010", 26071 => "00100011", 26073 => "01101011", 26075 => "00011010", 26076 => "11100000", 26079 => "01011000", 26080 => "01110000", 26081 => "01011000", 26082 => "01111111", 26083 => "10100100", 26084 => "11001001", 26085 => "00111111", 26087 => "00100111", 26088 => "01010100", 26095 => "00101101", 26099 => "01110010", 26100 => "01000110", 26101 => "10011101", 26102 => "01111010", 26103 => "01000100", 26106 => "01111001", 26110 => "00010100", 26111 => "11111010", 26113 => "10011101", 26115 => "10001010", 26116 => "11000111", 26117 => "11001101", 26118 => "10000011", 26119 => "01101100", 26120 => "11001011", 26124 => "01101101", 26127 => "11101100", 26129 => "10110001", 26130 => "01010010", 26135 => "11011010", 26136 => "11101001", 26138 => "10110111", 26139 => "00101000", 26142 => "00110001", 26143 => "00011001", 26144 => "11000001", 26145 => "10111111", 26147 => "01111011", 26149 => "01110101", 26153 => "11101101", 26156 => "10000010", 26158 => "11001111", 26159 => "01011111", 26160 => "01001111", 26163 => "11100100", 26165 => "10001010", 26166 => "10111001", 26167 => "01110111", 26169 => "01001101", 26170 => "01011100", 26171 => "11101110", 26172 => "01011001", 26174 => "11000011", 26177 => "10001010", 26178 => "10100000", 26185 => "10110011", 26187 => "00000110", 26188 => "10010100", 26189 => "01101101", 26191 => "10111001", 26193 => "11000110", 26194 => "11100101", 26195 => "11011100", 26196 => "10010000", 26197 => "11010000", 26202 => "00110110", 26203 => "10101110", 26204 => "00111110", 26205 => "00000111", 26208 => "00001011", 26210 => "10001000", 26217 => "01010001", 26218 => "01000010", 26219 => "00000110", 26222 => "11111100", 26223 => "10110100", 26224 => "00111111", 26225 => "01011010", 26230 => "10001111", 26235 => "01000001", 26236 => "01000111", 26238 => "11111110", 26241 => "11001011", 26242 => "10111111", 26243 => "11000011", 26245 => "01101101", 26248 => "10011100", 26249 => "01000110", 26254 => "00100011", 26255 => "10111000", 26256 => "11001100", 26257 => "10011110", 26259 => "11110110", 26260 => "01011101", 26261 => "11011001", 26263 => "11000111", 26265 => "00100010", 26266 => "10110101", 26270 => "01101010", 26272 => "01101101", 26273 => "10101011", 26276 => "00100000", 26279 => "11000111", 26280 => "11011011", 26283 => "00110010", 26285 => "00110010", 26287 => "10100010", 26288 => "11100010", 26290 => "11000011", 26293 => "10000011", 26294 => "00110101", 26296 => "01010001", 26297 => "11001110", 26298 => "11100010", 26300 => "01111010", 26301 => "00100010", 26303 => "11101010", 26304 => "01001110", 26307 => "01001110", 26308 => "01111100", 26309 => "00011111", 26311 => "11101010", 26312 => "11100011", 26314 => "10001011", 26315 => "11101111", 26317 => "00001101", 26319 => "10110011", 26320 => "11000100", 26322 => "11000111", 26324 => "01001011", 26326 => "11001011", 26328 => "00001111", 26329 => "00100000", 26333 => "01111010", 26334 => "11111001", 26335 => "00010110", 26336 => "10000100", 26337 => "10010011", 26338 => "01101001", 26339 => "01111010", 26341 => "01100011", 26344 => "01101011", 26347 => "10111000", 26350 => "10110100", 26352 => "11010111", 26353 => "00010110", 26354 => "01010110", 26355 => "01110111", 26356 => "10000101", 26361 => "10111100", 26362 => "01101010", 26363 => "10100010", 26364 => "10000110", 26365 => "10101011", 26366 => "10111010", 26367 => "01100010", 26368 => "11010110", 26372 => "01010011", 26374 => "10101100", 26375 => "01011011", 26379 => "10001110", 26380 => "11000100", 26381 => "10011011", 26382 => "00100110", 26388 => "00111001", 26392 => "10101101", 26393 => "11000000", 26394 => "10001111", 26395 => "11001010", 26396 => "00001011", 26397 => "00101011", 26398 => "10010011", 26400 => "11001000", 26401 => "10111011", 26403 => "11010101", 26404 => "10100000", 26407 => "11101101", 26413 => "00111110", 26416 => "00101001", 26417 => "11100111", 26419 => "10001000", 26425 => "10111101", 26428 => "11000110", 26429 => "10001001", 26435 => "11011100", 26436 => "00100110", 26437 => "00000011", 26438 => "11011010", 26439 => "00000001", 26440 => "00001111", 26443 => "00100101", 26447 => "01011110", 26448 => "11101001", 26450 => "10110101", 26451 => "00111111", 26452 => "00011010", 26458 => "10001111", 26460 => "11100010", 26461 => "11001010", 26467 => "11000000", 26469 => "00001100", 26470 => "00010011", 26471 => "00110001", 26472 => "01110001", 26473 => "01110001", 26475 => "11000011", 26476 => "10001011", 26480 => "11011010", 26481 => "11010000", 26484 => "00100011", 26485 => "00001000", 26486 => "00000001", 26487 => "10110000", 26490 => "00111001", 26491 => "00100001", 26492 => "10001100", 26495 => "11101010", 26497 => "11001110", 26498 => "10000101", 26499 => "11010010", 26500 => "10101011", 26501 => "11000100", 26502 => "01011011", 26503 => "00111011", 26505 => "11000111", 26507 => "00000111", 26510 => "11001100", 26511 => "10010011", 26513 => "11011111", 26514 => "11100101", 26515 => "01111010", 26516 => "01101001", 26517 => "00000010", 26518 => "01101101", 26519 => "00010100", 26523 => "10110000", 26524 => "00100100", 26525 => "00110110", 26528 => "10110010", 26529 => "01010110", 26530 => "01101100", 26532 => "00101101", 26537 => "11101000", 26549 => "00011110", 26551 => "00111111", 26554 => "11101101", 26557 => "00010100", 26559 => "00001111", 26562 => "10111110", 26564 => "11010010", 26567 => "00011001", 26568 => "10100011", 26569 => "11010101", 26573 => "11100011", 26574 => "00101101", 26575 => "01110001", 26577 => "01001101", 26579 => "11000001", 26580 => "10101100", 26581 => "10110010", 26582 => "11011111", 26584 => "10001111", 26586 => "10011000", 26587 => "01111101", 26590 => "01110010", 26594 => "01010111", 26599 => "10000111", 26600 => "11011000", 26601 => "10101111", 26604 => "10110110", 26605 => "01110001", 26607 => "01101110", 26609 => "10010001", 26611 => "10001111", 26612 => "11100010", 26614 => "00111111", 26615 => "00011001", 26617 => "00000110", 26620 => "11111011", 26622 => "00111010", 26625 => "10001011", 26627 => "00100110", 26631 => "01010111", 26633 => "11001100", 26634 => "10100010", 26635 => "11100010", 26640 => "11001111", 26641 => "10100111", 26643 => "11001010", 26648 => "11011110", 26649 => "11001011", 26650 => "01100010", 26651 => "10011101", 26652 => "10100010", 26654 => "01001111", 26662 => "11100000", 26664 => "01101100", 26667 => "11111010", 26668 => "00010010", 26670 => "01010000", 26671 => "00011010", 26672 => "11011010", 26673 => "00011011", 26675 => "11110001", 26676 => "01010000", 26678 => "11100101", 26679 => "00010101", 26683 => "01001101", 26684 => "10001100", 26685 => "10011110", 26687 => "01110100", 26688 => "00010101", 26691 => "00001001", 26692 => "01001000", 26698 => "11010110", 26699 => "11100100", 26701 => "11000000", 26703 => "01000011", 26705 => "11001000", 26708 => "01100110", 26710 => "01010101", 26715 => "01110101", 26716 => "10001110", 26717 => "11001000", 26718 => "11100100", 26719 => "01001001", 26720 => "11010110", 26721 => "00100010", 26722 => "10111000", 26723 => "11100000", 26725 => "11101101", 26727 => "01110011", 26728 => "01100110", 26729 => "00101001", 26730 => "00011110", 26734 => "10001010", 26736 => "11011011", 26743 => "01100101", 26746 => "11101100", 26747 => "10111010", 26751 => "00100101", 26752 => "10011110", 26753 => "00111110", 26754 => "10100101", 26755 => "11101101", 26756 => "00010011", 26759 => "11110101", 26760 => "10111100", 26763 => "11010011", 26764 => "00100111", 26765 => "00111001", 26766 => "01100101", 26767 => "01111010", 26768 => "10000101", 26770 => "10001011", 26772 => "10101110", 26773 => "11010100", 26774 => "00110101", 26775 => "01010110", 26778 => "00010101", 26780 => "11001000", 26781 => "10000110", 26783 => "00110010", 26784 => "10101110", 26785 => "10111111", 26786 => "01001011", 26788 => "00111101", 26789 => "01011101", 26790 => "01000010", 26791 => "01001010", 26792 => "11110111", 26795 => "11110011", 26796 => "01010011", 26797 => "01011011", 26798 => "11010100", 26799 => "11010000", 26800 => "11110110", 26802 => "01111010", 26803 => "10101100", 26804 => "10000111", 26806 => "01100100", 26807 => "11111110", 26809 => "01001110", 26811 => "10101011", 26812 => "00011010", 26814 => "01010110", 26817 => "10001100", 26822 => "01011100", 26823 => "00000110", 26824 => "11101001", 26825 => "10010001", 26826 => "00111011", 26827 => "11111000", 26829 => "01110000", 26832 => "11000010", 26835 => "11000010", 26837 => "11010001", 26838 => "01100001", 26839 => "10010010", 26840 => "00011010", 26841 => "10111111", 26844 => "11001111", 26845 => "00101000", 26846 => "10000000", 26848 => "00111001", 26850 => "11101111", 26851 => "00001111", 26852 => "11000110", 26853 => "00011101", 26858 => "10001100", 26859 => "00100100", 26861 => "10110110", 26864 => "00100000", 26866 => "00000110", 26870 => "10101010", 26871 => "10010010", 26875 => "11101010", 26876 => "00111010", 26877 => "11011100", 26879 => "00010010", 26884 => "11100100", 26885 => "00000101", 26886 => "01010001", 26889 => "10010101", 26890 => "11111001", 26891 => "11001111", 26892 => "11110001", 26893 => "11101011", 26894 => "00100110", 26895 => "01000011", 26896 => "10100100", 26897 => "10001000", 26898 => "00011100", 26899 => "00111100", 26900 => "00110100", 26901 => "01000010", 26904 => "11100001", 26907 => "10011101", 26908 => "10110010", 26913 => "00100100", 26915 => "01101100", 26919 => "11000011", 26920 => "11011110", 26922 => "11110011", 26923 => "01101111", 26929 => "00000011", 26931 => "00111110", 26934 => "11011110", 26935 => "00111001", 26937 => "11001010", 26943 => "00100100", 26946 => "00011111", 26947 => "01110110", 26948 => "01001010", 26950 => "01010000", 26958 => "00010010", 26959 => "10101111", 26960 => "10101110", 26966 => "11110100", 26967 => "00000110", 26970 => "00100010", 26973 => "10100010", 26974 => "10010100", 26976 => "11110011", 26977 => "01101101", 26979 => "00001101", 26981 => "00011010", 26983 => "01111001", 26984 => "10010101", 26987 => "00001111", 26988 => "00111100", 26989 => "01001011", 26992 => "01010011", 26997 => "11000110", 27001 => "00001111", 27002 => "01000011", 27003 => "11110100", 27005 => "11111111", 27006 => "00100000", 27008 => "01001010", 27012 => "10110101", 27013 => "01010110", 27024 => "10011100", 27025 => "11000110", 27026 => "00010001", 27029 => "01001111", 27032 => "11001111", 27036 => "11111100", 27037 => "00011101", 27038 => "00010001", 27039 => "11001100", 27041 => "00000100", 27042 => "11000101", 27044 => "00101011", 27045 => "00011101", 27046 => "11011111", 27047 => "01011000", 27050 => "00100100", 27052 => "01011011", 27056 => "10111000", 27059 => "01010110", 27060 => "01010111", 27063 => "00111011", 27065 => "10111101", 27070 => "10001111", 27073 => "00111101", 27075 => "00100000", 27084 => "11101101", 27085 => "00111000", 27086 => "11011101", 27088 => "10111011", 27090 => "00101111", 27093 => "01110010", 27094 => "01101001", 27095 => "11100011", 27098 => "10111111", 27102 => "01100110", 27104 => "11101110", 27105 => "11011010", 27107 => "11011010", 27112 => "11101111", 27113 => "11111110", 27114 => "11011101", 27117 => "10000101", 27118 => "11111011", 27120 => "00110010", 27121 => "00011001", 27122 => "01011111", 27124 => "10101010", 27126 => "01011100", 27128 => "11111110", 27129 => "00001100", 27130 => "11000010", 27132 => "10000010", 27133 => "11101100", 27136 => "00011011", 27141 => "11011011", 27144 => "11101101", 27145 => "00010001", 27148 => "11010011", 27152 => "00111110", 27153 => "00111001", 27157 => "11010011", 27158 => "01111100", 27159 => "01110110", 27168 => "10111011", 27173 => "01111111", 27174 => "10110100", 27177 => "11001001", 27180 => "10000101", 27182 => "10000110", 27183 => "00110101", 27184 => "00100100", 27187 => "10010001", 27188 => "00011111", 27191 => "11110011", 27192 => "00101001", 27195 => "00011111", 27197 => "10100100", 27200 => "01101110", 27203 => "01001110", 27206 => "00010001", 27209 => "01001101", 27210 => "11101010", 27211 => "10000110", 27215 => "01010101", 27217 => "10100011", 27218 => "01100010", 27220 => "11110010", 27221 => "10110100", 27222 => "01111000", 27223 => "00111101", 27225 => "10000101", 27229 => "00001001", 27231 => "11111100", 27233 => "10010010", 27234 => "10110100", 27236 => "10111111", 27237 => "00000010", 27245 => "10001100", 27247 => "10111010", 27249 => "11011101", 27252 => "10011000", 27253 => "01000101", 27254 => "01010111", 27258 => "10100010", 27259 => "00001010", 27262 => "01000000", 27264 => "01100110", 27265 => "10100110", 27267 => "11001110", 27268 => "00011111", 27269 => "01101011", 27270 => "00010101", 27271 => "01011110", 27274 => "01011000", 27275 => "01110010", 27281 => "00000101", 27282 => "01010010", 27283 => "10111111", 27288 => "11001101", 27290 => "10000111", 27291 => "11010111", 27292 => "00110011", 27293 => "10100011", 27294 => "00110000", 27295 => "01110111", 27298 => "11010111", 27301 => "10000001", 27304 => "00111110", 27306 => "01011111", 27307 => "00110110", 27309 => "01111111", 27310 => "01100110", 27312 => "10011000", 27313 => "00100010", 27315 => "10001011", 27316 => "01011110", 27317 => "01001101", 27322 => "01001110", 27325 => "10011001", 27326 => "11011100", 27328 => "01000001", 27330 => "00100100", 27332 => "10000001", 27333 => "10110001", 27336 => "10110001", 27338 => "10000010", 27341 => "01110011", 27345 => "01010101", 27348 => "00111011", 27349 => "10100100", 27350 => "11101101", 27351 => "10101001", 27352 => "01111001", 27354 => "01111001", 27355 => "01111100", 27358 => "00110001", 27362 => "11111110", 27363 => "11100111", 27365 => "01011000", 27369 => "01001001", 27372 => "00110111", 27373 => "10100001", 27376 => "00111111", 27380 => "11101100", 27381 => "10000011", 27382 => "00101000", 27385 => "00101110", 27387 => "00001100", 27388 => "10001010", 27389 => "00010000", 27390 => "10011000", 27391 => "11101100", 27392 => "11101101", 27393 => "11001001", 27395 => "11000011", 27396 => "01011000", 27398 => "11110101", 27400 => "10010001", 27401 => "11100101", 27406 => "01010010", 27407 => "11111000", 27408 => "10110011", 27409 => "10000001", 27410 => "10001011", 27412 => "11001111", 27417 => "10110101", 27418 => "00100000", 27419 => "10010111", 27421 => "00111001", 27423 => "01101101", 27424 => "01110011", 27429 => "01011100", 27433 => "01100111", 27435 => "10111010", 27438 => "10111000", 27440 => "11101010", 27441 => "01010010", 27443 => "01011111", 27444 => "10000110", 27445 => "10101011", 27446 => "00010111", 27449 => "00110001", 27450 => "00001100", 27451 => "00110001", 27452 => "11100000", 27454 => "11101101", 27455 => "00111010", 27458 => "10101111", 27459 => "00100110", 27460 => "01100011", 27461 => "10001101", 27464 => "11010111", 27465 => "10000101", 27466 => "00011101", 27468 => "11110010", 27470 => "10001110", 27471 => "01100111", 27474 => "01100001", 27475 => "10100011", 27478 => "01111001", 27479 => "00110011", 27480 => "11111001", 27481 => "10100101", 27483 => "10001100", 27486 => "11110111", 27487 => "10001101", 27488 => "11111000", 27489 => "00010001", 27490 => "11101100", 27491 => "00101011", 27493 => "01100110", 27495 => "10111001", 27496 => "11001100", 27498 => "11011100", 27500 => "01001100", 27507 => "10111001", 27510 => "00110101", 27511 => "10011101", 27512 => "11010000", 27514 => "01110110", 27516 => "00011010", 27517 => "01110000", 27519 => "11110000", 27522 => "00101000", 27524 => "00001001", 27527 => "01001101", 27530 => "11111010", 27531 => "10111010", 27533 => "11011101", 27534 => "01111111", 27536 => "10001011", 27541 => "00010101", 27542 => "10111001", 27543 => "01000001", 27545 => "11000110", 27546 => "01001000", 27547 => "00000010", 27549 => "01010110", 27551 => "00100000", 27553 => "00101111", 27555 => "10101001", 27559 => "01101101", 27560 => "00111000", 27562 => "00010110", 27563 => "10011100", 27570 => "01010101", 27571 => "01000010", 27572 => "01001111", 27573 => "10001110", 27575 => "10111110", 27577 => "11110100", 27579 => "11000010", 27580 => "11010111", 27582 => "10111011", 27591 => "00100010", 27594 => "01100001", 27596 => "01011111", 27600 => "10010101", 27601 => "00111101", 27604 => "11111110", 27605 => "00110011", 27606 => "11100011", 27607 => "01011101", 27608 => "11010111", 27612 => "10100011", 27622 => "10100010", 27623 => "10101011", 27624 => "00111111", 27625 => "10010010", 27628 => "10101100", 27629 => "00001000", 27630 => "10000000", 27633 => "00010001", 27634 => "10011010", 27635 => "11001101", 27637 => "11011101", 27638 => "00110100", 27640 => "11000101", 27641 => "00010101", 27655 => "01001100", 27656 => "00101011", 27657 => "10001111", 27659 => "10100000", 27660 => "10001100", 27667 => "10000000", 27668 => "01110100", 27670 => "01011110", 27671 => "10101100", 27672 => "10000100", 27675 => "11001010", 27676 => "10101010", 27677 => "10100011", 27679 => "10000101", 27682 => "01010110", 27687 => "10010111", 27688 => "10111110", 27689 => "10100101", 27690 => "11011010", 27692 => "10101110", 27696 => "11110100", 27697 => "11000111", 27699 => "01110000", 27701 => "00101011", 27702 => "00011000", 27704 => "10000100", 27706 => "01011110", 27708 => "10101111", 27710 => "10010100", 27714 => "10001001", 27715 => "00000101", 27717 => "11001101", 27719 => "11000001", 27720 => "11001100", 27721 => "00100101", 27723 => "01010000", 27725 => "11110111", 27726 => "00100011", 27730 => "00011111", 27731 => "10000100", 27732 => "10111111", 27734 => "10011111", 27736 => "00101101", 27737 => "10010100", 27743 => "00100101", 27744 => "10011101", 27745 => "11101001", 27746 => "01011111", 27749 => "10110011", 27750 => "10010011", 27753 => "10111010", 27754 => "11000101", 27755 => "10001101", 27756 => "10111001", 27757 => "01110001", 27760 => "01000110", 27761 => "11101001", 27762 => "10010111", 27763 => "01101100", 27764 => "11001110", 27765 => "00111010", 27766 => "10111011", 27767 => "00000101", 27768 => "10111111", 27769 => "11100010", 27770 => "00110001", 27772 => "11111001", 27773 => "00000100", 27775 => "11100011", 27779 => "10001111", 27782 => "00100111", 27785 => "10100001", 27786 => "01011100", 27787 => "00000010", 27788 => "10000001", 27794 => "00100011", 27795 => "11100010", 27796 => "01100010", 27799 => "11111111", 27800 => "10111001", 27808 => "10111111", 27810 => "11011010", 27811 => "01011110", 27815 => "01101100", 27817 => "00101100", 27819 => "01000110", 27825 => "00001111", 27829 => "01000001", 27830 => "10011100", 27832 => "01110000", 27833 => "10001010", 27834 => "00011100", 27835 => "01011100", 27838 => "11010111", 27840 => "11011001", 27844 => "11101111", 27848 => "10001110", 27849 => "01001000", 27850 => "11101110", 27853 => "00100000", 27855 => "11011000", 27857 => "10101010", 27858 => "01101101", 27859 => "11100001", 27865 => "00100001", 27866 => "01110001", 27868 => "11001001", 27870 => "10000100", 27872 => "01001110", 27875 => "10101111", 27876 => "01000101", 27877 => "01100101", 27878 => "11010010", 27881 => "10010001", 27882 => "10011000", 27885 => "10100010", 27887 => "10010001", 27888 => "00110111", 27898 => "10010101", 27900 => "01111000", 27903 => "11000111", 27904 => "01101000", 27909 => "00100111", 27911 => "11011101", 27913 => "01100100", 27914 => "11001111", 27916 => "00001110", 27917 => "00001000", 27918 => "01110011", 27919 => "11110111", 27921 => "10011110", 27922 => "01100000", 27926 => "00001010", 27930 => "10111110", 27933 => "10101000", 27936 => "11010111", 27938 => "10100110", 27940 => "10010101", 27946 => "10101011", 27950 => "11001101", 27952 => "00101001", 27953 => "01110000", 27954 => "01110100", 27955 => "00100000", 27957 => "10100100", 27958 => "01000000", 27960 => "11111111", 27963 => "11000111", 27964 => "01010000", 27966 => "01101111", 27967 => "11100011", 27971 => "01001011", 27972 => "11010101", 27974 => "00001010", 27980 => "10110001", 27981 => "11100100", 27982 => "11011110", 27983 => "11010010", 27986 => "10000111", 27987 => "01100001", 27990 => "01010100", 27991 => "11010100", 27992 => "01101010", 27995 => "11110101", 27997 => "01110000", 27998 => "01011001", 28002 => "10101011", 28003 => "00001010", 28010 => "10110000", 28011 => "00111010", 28013 => "11100110", 28014 => "11011000", 28015 => "11100010", 28016 => "10101101", 28020 => "11010011", 28023 => "11001111", 28024 => "00000110", 28029 => "00010101", 28030 => "00011000", 28032 => "01111010", 28033 => "00110111", 28036 => "00110011", 28039 => "00001011", 28040 => "01011111", 28044 => "01011100", 28046 => "00101100", 28049 => "00100111", 28052 => "01000100", 28053 => "01001001", 28054 => "00000101", 28056 => "11010011", 28059 => "01000000", 28061 => "11011001", 28069 => "00100111", 28071 => "10000100", 28073 => "11010010", 28075 => "01000010", 28080 => "10101101", 28082 => "00110000", 28083 => "01110000", 28085 => "11000001", 28087 => "11010000", 28088 => "11011010", 28089 => "10100010", 28090 => "01001101", 28092 => "00100011", 28094 => "00110010", 28098 => "01110011", 28100 => "00100101", 28104 => "10011111", 28105 => "11001010", 28109 => "11111011", 28115 => "11110111", 28121 => "00101100", 28123 => "01001111", 28124 => "01101011", 28129 => "11010101", 28131 => "01100101", 28133 => "11010110", 28134 => "01101111", 28135 => "11110110", 28139 => "11101000", 28140 => "10011110", 28141 => "10011000", 28142 => "00101110", 28146 => "11010110", 28148 => "11100001", 28150 => "10101101", 28151 => "00111010", 28154 => "00001001", 28155 => "11000001", 28158 => "00100101", 28160 => "11100110", 28161 => "10011111", 28162 => "10101100", 28163 => "01001110", 28165 => "10011111", 28167 => "10011010", 28168 => "11111111", 28172 => "10001111", 28173 => "00011001", 28176 => "11111010", 28177 => "11111111", 28179 => "11111000", 28180 => "10101001", 28181 => "00110110", 28183 => "11011100", 28185 => "00101001", 28186 => "00100100", 28188 => "01001000", 28189 => "11111000", 28190 => "00001101", 28192 => "11110100", 28194 => "00001111", 28197 => "11110110", 28198 => "11001010", 28200 => "01111000", 28203 => "10000001", 28205 => "00011111", 28207 => "01010110", 28211 => "11100010", 28213 => "01010001", 28214 => "01100010", 28216 => "11001111", 28217 => "01000110", 28219 => "01111000", 28221 => "01110000", 28222 => "01100100", 28223 => "00110101", 28238 => "00010100", 28242 => "11110100", 28243 => "10110101", 28248 => "10101101", 28249 => "00010101", 28250 => "01111111", 28252 => "10101111", 28253 => "00010100", 28256 => "11111000", 28260 => "11100100", 28261 => "01010110", 28262 => "10110110", 28263 => "11100011", 28264 => "10101010", 28265 => "11111111", 28272 => "11100010", 28273 => "00011110", 28276 => "11000111", 28278 => "01011000", 28280 => "10000011", 28281 => "10011110", 28286 => "00010011", 28287 => "01000001", 28289 => "01010001", 28290 => "00001000", 28292 => "11011011", 28293 => "01011101", 28294 => "01111101", 28295 => "10011000", 28297 => "10001010", 28299 => "11111111", 28301 => "01101001", 28302 => "01100100", 28303 => "11110001", 28308 => "00011110", 28309 => "01111011", 28310 => "10010111", 28312 => "11100101", 28314 => "01101011", 28316 => "10100110", 28317 => "11001000", 28318 => "11001011", 28320 => "01001110", 28323 => "10101101", 28334 => "01110001", 28336 => "10010111", 28338 => "10001001", 28339 => "10110111", 28340 => "00001100", 28342 => "00110000", 28344 => "10001100", 28345 => "01101111", 28347 => "10011110", 28348 => "10101011", 28349 => "01001001", 28350 => "00111010", 28351 => "01111010", 28352 => "01000010", 28359 => "00101111", 28361 => "00011001", 28362 => "01100100", 28364 => "10000111", 28366 => "11001101", 28367 => "11011010", 28370 => "10111110", 28372 => "10111010", 28374 => "10011100", 28375 => "00010000", 28378 => "10110010", 28382 => "01101101", 28383 => "11011110", 28387 => "00001011", 28388 => "10110110", 28390 => "01011001", 28393 => "01110100", 28396 => "00100010", 28397 => "00011011", 28398 => "10001110", 28399 => "01101101", 28400 => "00010101", 28401 => "10101000", 28402 => "00011010", 28406 => "01110000", 28407 => "11111010", 28408 => "11100001", 28410 => "00011111", 28411 => "10111011", 28413 => "11101001", 28416 => "10110011", 28417 => "01001100", 28418 => "11110010", 28419 => "11111011", 28420 => "01001001", 28423 => "10110000", 28425 => "00011001", 28426 => "00010110", 28431 => "10111110", 28432 => "10001000", 28435 => "00010111", 28439 => "00100111", 28442 => "00101110", 28443 => "00100000", 28445 => "10000100", 28447 => "00011001", 28448 => "01100010", 28455 => "10011111", 28457 => "00010010", 28458 => "00101000", 28460 => "10100001", 28461 => "10111101", 28465 => "10000000", 28466 => "10101110", 28468 => "01001001", 28469 => "11101111", 28470 => "00101010", 28471 => "11111111", 28472 => "00011100", 28473 => "11001001", 28474 => "00110111", 28476 => "10100010", 28480 => "01101111", 28482 => "01011110", 28488 => "11101000", 28489 => "11100011", 28490 => "10110111", 28493 => "10101110", 28500 => "10110101", 28501 => "10111011", 28506 => "00011111", 28508 => "01101110", 28509 => "11111000", 28510 => "10110011", 28513 => "01011100", 28517 => "10111101", 28518 => "11001101", 28519 => "10101011", 28521 => "00011000", 28522 => "00000101", 28523 => "01000111", 28525 => "00101101", 28528 => "10111110", 28529 => "11000010", 28534 => "00001001", 28537 => "01011101", 28538 => "00111000", 28539 => "00011010", 28540 => "01100101", 28541 => "01011100", 28547 => "00001011", 28549 => "10001100", 28552 => "01011010", 28553 => "01010110", 28557 => "01001000", 28562 => "11001101", 28563 => "00011011", 28565 => "10000000", 28566 => "01010000", 28567 => "00001011", 28568 => "10011010", 28569 => "11000100", 28570 => "10010000", 28571 => "01001011", 28575 => "01011101", 28576 => "11100110", 28577 => "00010110", 28583 => "00010000", 28584 => "10100011", 28586 => "10111011", 28589 => "01011010", 28590 => "00010011", 28594 => "01011100", 28596 => "01001100", 28607 => "01010000", 28609 => "10000100", 28610 => "11101100", 28616 => "10010110", 28619 => "11110010", 28620 => "10011011", 28621 => "10000100", 28623 => "00010000", 28627 => "01111000", 28629 => "00000010", 28632 => "10101110", 28635 => "01110100", 28636 => "01001001", 28638 => "01011111", 28640 => "01000010", 28641 => "10101011", 28642 => "11010011", 28643 => "01001011", 28648 => "11000001", 28649 => "10000000", 28651 => "10001100", 28654 => "00001111", 28655 => "11110011", 28656 => "11110101", 28657 => "01000001", 28658 => "00110011", 28661 => "10100110", 28662 => "10101101", 28663 => "11010111", 28664 => "00010110", 28665 => "10101110", 28670 => "00000010", 28671 => "00011111", 28673 => "00001000", 28674 => "11010100", 28675 => "01010111", 28677 => "00001000", 28678 => "01100110", 28679 => "10010111", 28680 => "10111000", 28681 => "00010100", 28683 => "00010100", 28685 => "10000111", 28686 => "11010100", 28687 => "00111100", 28688 => "10010101", 28689 => "00101100", 28691 => "10000010", 28696 => "01011110", 28698 => "01000100", 28703 => "01110011", 28705 => "00111011", 28707 => "01101000", 28709 => "01101111", 28711 => "10000100", 28714 => "11101111", 28715 => "00110001", 28717 => "00101011", 28719 => "10110010", 28720 => "01010011", 28723 => "00111010", 28726 => "00011110", 28729 => "00010001", 28731 => "11101111", 28732 => "11101001", 28733 => "11010000", 28734 => "01100010", 28741 => "00110000", 28744 => "01101000", 28746 => "00010110", 28747 => "11101100", 28749 => "01011000", 28750 => "00110110", 28753 => "01011000", 28758 => "01100010", 28759 => "01010000", 28765 => "00100110", 28773 => "01000001", 28774 => "10111100", 28775 => "10111101", 28777 => "10111001", 28781 => "10110001", 28783 => "01100111", 28785 => "11110111", 28786 => "01000100", 28788 => "00001110", 28789 => "10000110", 28793 => "00010000", 28794 => "10001100", 28799 => "11100011", 28801 => "10001011", 28803 => "00100001", 28804 => "01100101", 28813 => "10110101", 28815 => "00101000", 28816 => "10100111", 28820 => "01100010", 28822 => "00110010", 28823 => "10111110", 28825 => "01110000", 28826 => "11001011", 28827 => "00101000", 28830 => "11000000", 28833 => "00000001", 28836 => "11001110", 28837 => "11101100", 28838 => "10000111", 28839 => "11001101", 28842 => "01010101", 28843 => "01101011", 28845 => "01010101", 28849 => "11110111", 28850 => "00011000", 28851 => "11011111", 28852 => "11000010", 28854 => "00011101", 28855 => "00111000", 28856 => "01010100", 28857 => "10001100", 28858 => "11111001", 28859 => "01110001", 28861 => "11000111", 28865 => "01010011", 28866 => "11111010", 28868 => "00101101", 28870 => "11011111", 28871 => "00101010", 28872 => "01011010", 28873 => "10100100", 28874 => "11000010", 28877 => "11010100", 28879 => "00111000", 28881 => "01011111", 28882 => "01100110", 28886 => "01100010", 28887 => "00110010", 28889 => "11100111", 28891 => "01100100", 28893 => "01011010", 28897 => "10110010", 28898 => "01001011", 28899 => "01110101", 28900 => "10001111", 28901 => "10000011", 28902 => "10011010", 28904 => "00001101", 28911 => "11111111", 28913 => "11111110", 28916 => "01000111", 28917 => "01110000", 28918 => "00111100", 28920 => "00110000", 28923 => "10110111", 28924 => "01011011", 28925 => "01001001", 28926 => "00000010", 28929 => "01100000", 28931 => "10011001", 28935 => "11010111", 28936 => "00100110", 28937 => "00011010", 28938 => "00100101", 28939 => "10001001", 28940 => "01011100", 28942 => "10101001", 28943 => "10101001", 28944 => "11001010", 28946 => "01100111", 28948 => "01001101", 28952 => "01111010", 28953 => "11010100", 28954 => "11011101", 28957 => "10101111", 28960 => "11000100", 28961 => "11101011", 28963 => "10110100", 28966 => "00001101", 28967 => "10100011", 28968 => "00100011", 28969 => "01111000", 28972 => "10100011", 28974 => "01110110", 28976 => "11000000", 28979 => "01111100", 28980 => "00100111", 28982 => "01010000", 28985 => "11100111", 28986 => "00100011", 28989 => "11010001", 28990 => "00000011", 28991 => "10000111", 28992 => "11110000", 28994 => "11010001", 28995 => "01011111", 28998 => "01111100", 29000 => "01010101", 29008 => "01010101", 29009 => "00000110", 29010 => "00110001", 29015 => "11100111", 29017 => "11110000", 29020 => "00101000", 29024 => "11011010", 29026 => "10000010", 29031 => "10100011", 29032 => "10000100", 29033 => "10011001", 29034 => "01000111", 29035 => "00001010", 29038 => "10111111", 29039 => "11001001", 29040 => "01100111", 29042 => "10001101", 29044 => "01001100", 29046 => "00001011", 29048 => "01010000", 29050 => "11101110", 29052 => "01101111", 29053 => "00001100", 29057 => "11011000", 29059 => "01010000", 29061 => "00011010", 29062 => "11010010", 29063 => "00011010", 29064 => "11001101", 29073 => "11110010", 29075 => "01000110", 29077 => "01011011", 29079 => "10101101", 29080 => "11101001", 29081 => "00001110", 29082 => "11010011", 29090 => "00111110", 29091 => "01110101", 29095 => "11110010", 29102 => "11011001", 29105 => "10100110", 29106 => "00011011", 29107 => "00000001", 29112 => "00001101", 29113 => "00111111", 29119 => "00100011", 29120 => "11001000", 29122 => "01110001", 29125 => "10000010", 29133 => "11011110", 29134 => "01011100", 29136 => "10111101", 29137 => "01010011", 29139 => "01001110", 29141 => "01011100", 29148 => "01011000", 29149 => "00001101", 29151 => "11101110", 29152 => "11011111", 29154 => "10001101", 29157 => "00101010", 29158 => "01100111", 29159 => "00110000", 29162 => "00100000", 29165 => "10100010", 29168 => "01001011", 29175 => "10100110", 29176 => "11100011", 29178 => "01011110", 29179 => "10111010", 29180 => "10100010", 29185 => "10111011", 29189 => "00011100", 29191 => "11110111", 29194 => "10101000", 29195 => "11001111", 29196 => "00001000", 29198 => "00010111", 29201 => "01110000", 29203 => "01001000", 29204 => "11001010", 29206 => "01000110", 29208 => "10011100", 29209 => "10011001", 29212 => "01010000", 29214 => "00110111", 29215 => "10110011", others => (others =>'0'));component project_reti_logiche is 
    port (
            i_clk         : in  std_logic;
            i_start       : in  std_logic;
            i_rst         : in  std_logic;
            i_data       : in  std_logic_vector(7 downto 0); --1 byte
            o_address     : out std_logic_vector(15 downto 0); --16 bit addr: max size is 255*255 + 3 more for max x and y and thresh.
            o_done            : out std_logic;
            o_en         : out std_logic;
            o_we       : out std_logic;
            o_data            : out std_logic_vector (7 downto 0)
          );
end component project_reti_logiche;


begin 
	UUT: project_reti_logiche
	port map (
		  i_clk      	=> tb_clk,	
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address, 
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
		  o_we 	=> mem_we,
          o_data    => mem_i_data
);

p_CLK_GEN : process is
  begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
  end process p_CLK_GEN; 
  
  
MEM : process(tb_clk)
   begin
    if tb_clk'event and tb_clk = '1' then
     if enable_wire = '1' then
      if mem_we = '1' then
       RAM(conv_integer(mem_address))              <= mem_i_data;
       mem_o_data                      <= mem_i_data after 1 ns;
      else
       mem_o_data <= RAM(conv_integer(mem_address)) after 1 ns;
      end if;
     end if;
    end if;
   end process;
 
  
test : process is
begin 
wait for 100 ns;
wait for c_CLOCK_PERIOD;
tb_rst <= '1';
wait for c_CLOCK_PERIOD;
tb_rst <= '0';
wait for c_CLOCK_PERIOD;
tb_start <= '1';
wait for c_CLOCK_PERIOD; 
tb_start <= '0';
wait until tb_done = '1';
wait until tb_done = '0';
wait until rising_edge(tb_clk); 

assert RAM(1) = "01110010" report "FAIL high bits" severity failure;
assert RAM(0) = "00100000" report "FAIL low bits" severity failure;
assert false report "Simulation Ended!, test passed" severity failure;
end process test;
end projecttb;