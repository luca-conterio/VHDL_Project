----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 12.12.2017 17:48:44
-- Design Name: 
-- Module Name: FSM_testbench - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
 
entity project_tb is
end project_tb;


architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 15 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst		    : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		    : std_logic := '0';
signal   mem_o_data,mem_i_data		: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		: std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (2 => "00010011", 3 => "00011110", 4 => "00000000", 7 => "01101011", 8 => "10011000", 11 => "01111010", 14 => "10001100", 17 => "11011110", 18 => "00001110", 19 => "01111100", 21 => "00111011", 24 => "10010100", 31 => "00000101", 34 => "01010001", 35 => "10000101", 36 => "00101001", 39 => "11000010", 40 => "01101111", 43 => "01010110", 44 => "11100100", 46 => "01011101", 50 => "11010110", 52 => "10011000", 54 => "10010100", 55 => "00001110", 57 => "10010100", 58 => "11010000", 59 => "11111011", 64 => "10011010", 65 => "10000110", 68 => "11011110", 76 => "11011110", 77 => "00000011", 78 => "11010001", 83 => "01111001", 84 => "00000111", 85 => "00100101", 87 => "11011011", 88 => "11110100", 89 => "10101100", 90 => "01011110", 92 => "01111001", 94 => "11101011", 96 => "01111010", 98 => "01010011", 100 => "11100101", 102 => "11111011", 103 => "11011101", 105 => "01001111", 108 => "11111100", 109 => "00110010", 111 => "11010111", 115 => "01001011", 117 => "11000100", 118 => "10110011", 119 => "01111101", 123 => "00000011", 125 => "00001001", 126 => "10110100", 127 => "00110010", 128 => "10001101", 134 => "11010000", 135 => "00001001", 136 => "11100101", 137 => "11010111", 139 => "10001100", 140 => "10011111", 142 => "00100010", 143 => "00110111", 147 => "01100110", 148 => "01111100", 149 => "01110101", 150 => "11011101", 153 => "11101110", 155 => "00000001", 160 => "00010110", 161 => "11111111", 172 => "10110001", 173 => "01110001", 174 => "00010101", 175 => "00111100", 177 => "00110110", 180 => "00001001", 181 => "01010010", 185 => "00000011", 186 => "01000101", 190 => "00010111", 191 => "00111100", 192 => "10110001", 194 => "00111110", 195 => "01011000", 198 => "11110011", 199 => "11011010", 201 => "11000111", 202 => "01111111", 205 => "01011101", 206 => "11111011", 207 => "10101100", 213 => "11001011", 214 => "01010101", 215 => "00110100", 216 => "01101100", 217 => "00001001", 219 => "10111001", 222 => "01010110", 223 => "01011100", 225 => "00000011", 226 => "01101000", 228 => "01001000", 230 => "10011100", 232 => "11000000", 233 => "00111000", 236 => "00110010", 237 => "10001000", 239 => "01100110", 241 => "10100010", 243 => "01000101", 247 => "10010100", 253 => "01010010", 254 => "11100000", 255 => "10011011", 256 => "11001010", 259 => "01011000", 260 => "01010010", 262 => "00110101", 264 => "10001010", 265 => "11111110", 266 => "11011111", 270 => "11001100", 272 => "01001110", 274 => "00101010", 275 => "01100101", 276 => "01001100", 278 => "11100101", 281 => "10111100", 282 => "00000100", 285 => "10001000", 286 => "10101010", 287 => "10000111", 288 => "01001100", 291 => "01001111", 295 => "00011101", 296 => "10000010", 298 => "01100001", 299 => "00000110", 305 => "01110110", 311 => "01111111", 312 => "01001111", 313 => "01001010", 314 => "00000111", 317 => "11101100", 318 => "11011111", 320 => "11000010", 321 => "00100101", 322 => "10010111", 323 => "10010010", 324 => "10011011", 325 => "11101000", 326 => "11000101", 328 => "00101110", 330 => "11110101", 331 => "11100000", 332 => "10010010", 333 => "00100000", 334 => "11001100", 335 => "11111010", 336 => "01110101", 338 => "00111110", 341 => "11001111", 342 => "11110011", 344 => "00110111", 346 => "10111001", 349 => "10110101", 352 => "10001010", 353 => "10100010", 355 => "01111001", 356 => "11111010", 358 => "01011011", 359 => "11111001", 361 => "10111000", 362 => "01001011", 366 => "11000110", 369 => "01100011", 370 => "00110010", 374 => "11001101", 376 => "10110111", 378 => "01101101", 379 => "11000101", 380 => "10101001", 381 => "01101010", 382 => "11000010", 384 => "00101000", 387 => "01101100", 396 => "10101010", 398 => "01100110", 400 => "10011001", 402 => "00011011", 403 => "00011010", 405 => "11011101", 407 => "11001101", 410 => "01110000", 414 => "01100101", 416 => "00100011", 419 => "11100011", 420 => "01100110", 423 => "01100001", 426 => "11110001", 429 => "11100110", 431 => "00000010", 433 => "00110010", 435 => "10100101", 436 => "01010100", 439 => "10001010", 440 => "11111110", 445 => "11101010", 446 => "01100001", 447 => "00001101", 448 => "01010110", 453 => "10010101", 454 => "10110011", 455 => "11000101", 460 => "01011010", 461 => "10001011", 462 => "01100001", 464 => "01011000", 466 => "10011001", 467 => "01110000", 473 => "00010010", 474 => "01001101", 480 => "01101110", 481 => "11000001", 483 => "01010010", 484 => "10111001", 487 => "01100010", 488 => "10100111", 490 => "10100100", 491 => "10111001", 492 => "01100110", 496 => "11110001", 500 => "01010010", 501 => "00011101", 503 => "10010110", 507 => "01001111", 508 => "10010101", 512 => "01000001", 515 => "00100100", 520 => "10001111", 521 => "00000011", 529 => "11011110", 530 => "10011100", 532 => "10111100", 533 => "10100110", 537 => "10000111", 538 => "10101011", 539 => "01010111", 540 => "00100010", 541 => "11101010", 542 => "11001010", 543 => "01111111", 544 => "00100001", 549 => "11101011", 550 => "10010111", 552 => "11011110", 553 => "11001101", 557 => "10011010", 560 => "10111001", 561 => "10011001", 562 => "11111100", 563 => "00101111", 564 => "10010111", 565 => "01010000", others => (others =>'0'));component project_reti_logiche is 
    port (
            i_clk         : in  std_logic;
            i_start       : in  std_logic;
            i_rst         : in  std_logic;
            i_data       : in  std_logic_vector(7 downto 0); --1 byte
            o_address     : out std_logic_vector(15 downto 0); --16 bit addr: max size is 255*255 + 3 more for max x and y and thresh.
            o_done            : out std_logic;
            o_en         : out std_logic;
            o_we       : out std_logic;
            o_data            : out std_logic_vector (7 downto 0)
          );
end component project_reti_logiche;


begin 
	UUT: project_reti_logiche
	port map (
		  i_clk      	=> tb_clk,	
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address, 
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
		  o_we 	=> mem_we,
          o_data    => mem_i_data
);

p_CLK_GEN : process is
  begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
  end process p_CLK_GEN; 
  
  
MEM : process(tb_clk)
   begin
    if tb_clk'event and tb_clk = '1' then
     if enable_wire = '1' then
      if mem_we = '1' then
       RAM(conv_integer(mem_address))              <= mem_i_data;
       mem_o_data                      <= mem_i_data after 1 ns;
      else
       mem_o_data <= RAM(conv_integer(mem_address)) after 1 ns;
      end if;
     end if;
    end if;
   end process;
 
  
test : process is
begin 
wait for 100 ns;
wait for c_CLOCK_PERIOD;
tb_rst <= '1';
wait for c_CLOCK_PERIOD;
tb_rst <= '0';
wait for c_CLOCK_PERIOD;
tb_start <= '1';
wait for c_CLOCK_PERIOD; 
tb_start <= '0';
wait until tb_done = '1';
wait until tb_done = '0';
wait until rising_edge(tb_clk); 

assert RAM(1) = "00000010" report "FAIL high bits" severity failure;
assert RAM(0) = "00111010" report "FAIL low bits" severity failure;
assert false report "Simulation Ended!, test passed" severity failure;
end process test;
end projecttb;