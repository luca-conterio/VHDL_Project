----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 12.12.2017 17:48:44
-- Design Name: 
-- Module Name: FSM_testbench - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
 
entity project_tb is
end project_tb;


architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 15 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst		    : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		    : std_logic := '0';
signal   mem_o_data,mem_i_data		: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		: std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (2 => "01110101", 3 => "11100110", 4 => "10100110", 5 => "10110100", 6 => "10011101", 7 => "00011110", 8 => "00000010", 10 => "10000000", 11 => "10111010", 12 => "00011111", 15 => "11010000", 16 => "10101111", 17 => "00100111", 19 => "01100000", 22 => "10010100", 23 => "00111110", 24 => "00101010", 25 => "11101001", 27 => "10101000", 28 => "11001011", 29 => "10100110", 30 => "01101101", 31 => "11000111", 32 => "11011010", 35 => "00101000", 37 => "00101001", 38 => "10011100", 39 => "00011100", 40 => "00010000", 41 => "10010010", 43 => "10011110", 46 => "00001001", 47 => "01001100", 48 => "11011101", 49 => "00011110", 50 => "01101011", 51 => "01000000", 52 => "00001010", 53 => "00101001", 54 => "11111011", 58 => "01010011", 59 => "01110101", 63 => "11011000", 64 => "10110000", 66 => "01010000", 67 => "10011011", 68 => "01111000", 69 => "01100100", 70 => "00111111", 71 => "01110010", 72 => "01000100", 73 => "10100011", 75 => "01101100", 76 => "10111001", 77 => "10100101", 78 => "11010010", 79 => "10101000", 81 => "00001101", 82 => "01100111", 83 => "00001011", 84 => "10000011", 87 => "11000011", 89 => "11001100", 90 => "10011101", 93 => "00110111", 94 => "00101000", 95 => "11000011", 96 => "00011001", 97 => "00011010", 100 => "10111011", 101 => "10011011", 103 => "00111001", 104 => "10100101", 106 => "10001110", 107 => "01011010", 110 => "00001100", 111 => "10011101", 112 => "00110111", 113 => "11111100", 115 => "11101111", 116 => "11101101", 119 => "11101011", 120 => "00101010", 121 => "00011011", 122 => "11000001", 123 => "11110101", 124 => "11110001", 125 => "11000010", 127 => "10101011", 128 => "10111000", 129 => "10000100", 133 => "00010100", 134 => "00100111", 135 => "11101110", 136 => "10010011", 137 => "01010110", 138 => "00010101", 139 => "10111110", 142 => "11001101", 143 => "11010101", 144 => "01001111", 145 => "11110100", 146 => "11010001", 147 => "00010100", 148 => "01000000", 149 => "10000110", 150 => "11101011", 151 => "01010001", 152 => "10101101", 153 => "11011011", 154 => "00010000", 155 => "00111000", 156 => "00100010", 157 => "11000000", 158 => "00010010", 161 => "11001100", 162 => "00010100", 164 => "10011100", 166 => "11000111", 167 => "10101110", 168 => "10110011", 170 => "11011011", 171 => "00001111", 173 => "11011101", 174 => "00011010", 175 => "11001000", 176 => "11110010", 177 => "00010010", 178 => "00111101", 179 => "10111111", 180 => "01110111", 182 => "11010010", 183 => "10110010", 184 => "10111100", 185 => "11110100", 187 => "11100100", 188 => "11001100", 190 => "00001111", 191 => "00111000", 192 => "10010111", 193 => "00100000", 194 => "00100000", 195 => "11001000", 196 => "10111000", 197 => "00111111", 198 => "10010010", 199 => "10011001", 201 => "00010010", 202 => "11111110", 203 => "10110101", 204 => "10010100", 205 => "10000000", 206 => "11001011", 207 => "10100000", 208 => "00011000", 209 => "11011011", 210 => "00100110", 212 => "11111101", 214 => "00001101", 215 => "00111010", 216 => "00101000", 217 => "00000010", 218 => "00100001", 219 => "00010110", 220 => "11010101", 221 => "11111110", 222 => "10111000", 224 => "00110111", 225 => "01110111", 227 => "11111100", 228 => "00100000", 231 => "11010000", 232 => "10111111", 233 => "00010100", 235 => "01110101", 236 => "00101001", 237 => "11110101", 238 => "01000000", 239 => "00110111", 240 => "01111010", 241 => "10101110", 242 => "01101011", 243 => "00100010", 246 => "10101011", 248 => "01000111", 249 => "10001100", 250 => "00110011", 251 => "01101110", 254 => "11011100", 255 => "00011111", 258 => "01010110", 259 => "10000010", 260 => "11101100", 263 => "01000100", 264 => "01111101", 265 => "10111000", 266 => "10011010", 268 => "10110011", 269 => "01001011", 271 => "11001001", 272 => "11110000", 274 => "01101001", 277 => "00111101", 278 => "11001111", 280 => "10110111", 281 => "11110100", 282 => "10101110", 284 => "10101001", 288 => "00111110", 289 => "11000011", 291 => "01101111", 293 => "10010111", 294 => "00001010", 295 => "00100100", 296 => "10100100", 298 => "10011010", 302 => "00010010", 303 => "00100101", 304 => "10000110", 306 => "00000110", 307 => "11111001", 308 => "11010010", 309 => "11000100", 310 => "00000001", 311 => "01110110", 312 => "00001111", 313 => "10000000", 315 => "01000110", 316 => "11011100", 317 => "01100001", 319 => "10010110", 320 => "01101100", 321 => "10010100", 322 => "11101110", 324 => "00101110", 326 => "00101101", 327 => "00010100", 329 => "10111101", 330 => "10001010", 331 => "10000111", 332 => "11111000", 333 => "11111111", 334 => "11011000", 336 => "11000011", 337 => "10100000", 338 => "11001100", 339 => "01110111", 341 => "01100101", 342 => "01110010", 343 => "00010010", 344 => "01010001", 346 => "00100101", 347 => "01000011", 349 => "10100101", 351 => "00001010", 352 => "11010101", 353 => "00001000", 354 => "00101010", 355 => "00100111", 356 => "01011000", 357 => "00011101", 359 => "10100000", 361 => "01110111", 363 => "10100001", 365 => "11011011", 366 => "11100101", 367 => "10110001", 368 => "11000111", 369 => "11111011", 370 => "01110110", 371 => "01000010", 372 => "11101001", 373 => "01010010", 375 => "11100011", 377 => "00101100", 378 => "11100110", 379 => "10000000", 381 => "00011100", 383 => "10111001", 384 => "01001100", 385 => "11101101", 386 => "11000000", 387 => "01101110", 389 => "01101100", 390 => "11011110", 391 => "11101011", 392 => "10011100", 395 => "11101011", 396 => "11101111", 397 => "00100101", 398 => "01000011", 400 => "00001011", 401 => "10111101", 404 => "01101011", 406 => "10111011", 407 => "10101100", 408 => "10100001", 409 => "00011101", 410 => "00110011", 411 => "00111111", 413 => "00000101", 414 => "10011010", 415 => "01000010", 416 => "01110000", 418 => "01000110", 419 => "00010001", 421 => "10011111", 424 => "10010100", 426 => "10011001", 427 => "11010100", 428 => "10111100", 429 => "10111001", 430 => "01101100", 431 => "11111000", 433 => "01010100", 434 => "10010101", 435 => "10100110", 436 => "01100100", 437 => "11001110", 438 => "01110111", 439 => "10101100", 441 => "00100000", 442 => "10001101", 443 => "10011111", 444 => "01101011", 446 => "00011000", 447 => "10110101", 449 => "11010111", 450 => "01101010", 451 => "10111000", 452 => "10010101", 454 => "00100101", 455 => "00110111", 456 => "00101111", 457 => "10001000", 458 => "10110000", 459 => "10010100", 461 => "01010011", 462 => "11101000", 465 => "01100000", 466 => "11101100", 467 => "01100111", 468 => "00001101", 469 => "10111001", 470 => "11111101", 471 => "10111011", 472 => "10100111", 473 => "01100100", 475 => "01110010", 476 => "10101000", 477 => "10100011", 480 => "10011000", 481 => "11011110", 482 => "10100000", 483 => "10001101", 484 => "11010000", 486 => "11011111", 488 => "01111111", 490 => "11011111", 491 => "11110100", 492 => "11101101", 493 => "10011000", 494 => "10110001", 495 => "00001011", 496 => "01011011", 497 => "11100011", 499 => "10000000", 502 => "00011011", 503 => "01011110", 504 => "10010100", 505 => "01001011", 506 => "10110010", 507 => "10111111", 510 => "11011010", 511 => "01111010", 512 => "00111111", 513 => "10000011", 514 => "00001101", 515 => "01010010", 516 => "11000000", 517 => "10110101", 518 => "00111010", 519 => "10100111", 520 => "01010100", 521 => "11001111", 522 => "10111000", 524 => "00011101", 525 => "00010100", 527 => "11001000", 528 => "01101000", 529 => "11111100", 530 => "10010000", 531 => "01111101", 532 => "11111110", 533 => "00101001", 536 => "01011101", 537 => "00011011", 539 => "01010001", 540 => "00000100", 541 => "00101101", 542 => "10111011", 543 => "11000001", 549 => "11101110", 550 => "00000100", 553 => "11100011", 554 => "01010101", 555 => "01111100", 556 => "01001110", 557 => "01110010", 560 => "10001110", 561 => "00001110", 562 => "10011100", 563 => "01110010", 564 => "11010100", 566 => "01001110", 567 => "00110111", 570 => "01100100", 571 => "10010001", 572 => "00111101", 573 => "11101101", 574 => "10000100", 575 => "00100001", 576 => "00010101", 578 => "00101000", 579 => "00010000", 581 => "00000100", 583 => "11001100", 585 => "00011011", 586 => "00110001", 587 => "00001101", 589 => "00011100", 590 => "01111111", 591 => "10101001", 592 => "01010001", 593 => "00001000", 594 => "11011101", 595 => "11111101", 596 => "11011110", 597 => "11001101", 599 => "00100000", 600 => "11111110", 601 => "10101111", 602 => "10110111", 603 => "10000110", 604 => "01000010", 606 => "00111011", 607 => "11111100", 611 => "01001100", 612 => "00001000", 613 => "11010011", 614 => "01001001", 615 => "01100001", 616 => "10110100", 617 => "00111001", 618 => "11001100", 620 => "10001000", 623 => "01011001", 624 => "10011000", 625 => "11001101", 627 => "10110010", 630 => "11100111", 632 => "11011111", 633 => "11101001", 634 => "01010001", 636 => "00111101", 637 => "00010001", 640 => "01101101", 641 => "00001000", 642 => "01111010", 643 => "01000001", 644 => "10010001", 645 => "00010110", 647 => "01110111", 648 => "01111000", 649 => "10111111", 650 => "11010000", 651 => "01010011", 652 => "10001110", 654 => "10010100", 655 => "11011000", 656 => "01111010", 657 => "00110100", 658 => "10101000", 660 => "00010010", 662 => "01010110", 664 => "11100010", 665 => "10010110", 666 => "10011111", 667 => "11000101", 668 => "01111110", 670 => "01001011", 671 => "11010010", 672 => "11010100", 674 => "01111011", 675 => "11001000", 677 => "01001110", 678 => "00110101", 679 => "11101110", 680 => "11010101", 681 => "11100101", 683 => "10000111", 684 => "11001110", 685 => "10101110", 686 => "01010010", 687 => "00011001", 688 => "01100111", 689 => "01111101", 691 => "10101110", 692 => "01011110", 693 => "10011011", 694 => "01110110", 695 => "10100011", 698 => "00001111", 701 => "10101100", 702 => "11010011", 703 => "01100010", 704 => "11011101", 706 => "11000101", 707 => "11001111", 708 => "11001010", 709 => "01010011", 710 => "10011110", 711 => "01100100", 713 => "10111011", 716 => "11101100", 717 => "01000001", 718 => "01000110", 721 => "00011100", 724 => "00010100", 725 => "11100000", 728 => "11011011", 729 => "10110001", 730 => "11000111", 731 => "01110101", 734 => "11011011", 735 => "10101001", 736 => "00001100", 737 => "00100000", 741 => "01010100", 742 => "01011100", 743 => "11011101", 744 => "11100000", 746 => "11000101", 748 => "01000101", 750 => "10001100", 751 => "00101010", 752 => "00110110", 753 => "11001011", 754 => "11000000", 755 => "00101111", 756 => "00000100", 758 => "01010111", 759 => "01000101", 761 => "01101110", 762 => "10100000", 765 => "01100000", 767 => "11111000", 768 => "01000110", 771 => "11101101", 772 => "10010111", 773 => "10111001", 774 => "10101100", 775 => "11111000", 777 => "01001100", 780 => "00010100", 781 => "11010101", 782 => "01100100", 783 => "10001010", 784 => "10110100", 785 => "00101100", 786 => "01110000", 787 => "10111011", 788 => "10110111", 789 => "11100110", 790 => "01000001", 792 => "00111100", 793 => "10100010", 794 => "10011010", 796 => "01001111", 799 => "11010000", 801 => "11011000", 802 => "11101101", 805 => "01110111", 806 => "01100001", 808 => "00100111", 809 => "11110110", 810 => "10011101", 811 => "00100011", 812 => "00110011", 813 => "00111100", 815 => "00010101", 816 => "10101110", 817 => "01110100", 818 => "10111000", 822 => "00001011", 823 => "01111001", 826 => "01110111", 828 => "10110100", 829 => "01110110", 830 => "01000110", 834 => "00101101", 835 => "01000011", 836 => "10111100", 837 => "10110010", 838 => "11011010", 839 => "01101110", 840 => "01011001", 841 => "01101000", 844 => "01000001", 845 => "00100101", 846 => "00011001", 847 => "00000110", 848 => "11111100", 849 => "00100101", 850 => "10110011", 852 => "01000000", 853 => "10000011", 854 => "10000101", 856 => "01000000", 857 => "00000111", 860 => "01000001", 861 => "11100000", 863 => "00011011", 864 => "00101101", 865 => "10110001", 867 => "11111100", 868 => "10110110", 870 => "01011111", 872 => "11100100", 874 => "00101000", 875 => "00011000", 876 => "00010111", 877 => "11000010", 878 => "11110111", 881 => "10100100", 882 => "01110100", 886 => "00110110", 887 => "11100110", 888 => "01000111", 889 => "10010001", 890 => "11100100", 891 => "10101010", 892 => "01000110", 893 => "11110111", 894 => "00110001", 896 => "11101011", 897 => "11101001", 898 => "01001101", 899 => "00010100", 900 => "11011100", 901 => "01010000", 902 => "00000100", 903 => "01001111", 905 => "11100010", 906 => "00110110", 907 => "10100111", 908 => "01011101", 912 => "11111110", 913 => "10111110", 914 => "00001101", 915 => "00101101", 917 => "10001101", 919 => "11100000", 920 => "00000100", 921 => "00110110", 922 => "01010010", 923 => "01111101", 924 => "11101000", 925 => "10011100", 926 => "00010011", 927 => "11110011", 928 => "11101001", 929 => "01011011", 930 => "01000110", 933 => "10010111", 935 => "01010110", 937 => "00111110", 938 => "01100011", 941 => "11111101", 943 => "00001001", 945 => "01101110", 946 => "10010010", 948 => "11100001", 950 => "00010011", 951 => "00011110", 954 => "01001111", 956 => "11001111", 957 => "10011000", 958 => "00100111", 960 => "11001100", 963 => "10000010", 964 => "10110101", 966 => "10111100", 967 => "10100011", 968 => "00000001", 969 => "01110000", 972 => "10111000", 974 => "01011111", 975 => "01011110", 977 => "00011001", 978 => "01100011", 979 => "11010011", 980 => "01000101", 981 => "01110000", 985 => "00111100", 986 => "00111110", 987 => "10010110", 988 => "11110000", 989 => "00110100", 990 => "11010100", 991 => "10011100", 993 => "11010001", 994 => "01010100", 995 => "01101111", 998 => "11110010", 1000 => "00101011", 1001 => "10110000", 1003 => "01110111", 1004 => "00111111", 1007 => "10000110", 1008 => "00011110", 1009 => "10101100", 1010 => "00010101", 1011 => "10110111", 1012 => "11010100", 1013 => "11011001", 1015 => "01111000", 1017 => "10001010", 1018 => "00110110", 1019 => "01000000", 1020 => "00101001", 1021 => "10110010", 1022 => "01010111", 1023 => "10111111", 1024 => "01000000", 1027 => "10010100", 1028 => "01110010", 1030 => "11011111", 1031 => "00100111", 1033 => "01101011", 1034 => "11111011", 1035 => "00100101", 1036 => "10111110", 1037 => "00011101", 1038 => "01011001", 1040 => "01000111", 1041 => "11100000", 1042 => "00001010", 1043 => "00001011", 1044 => "01101011", 1045 => "00000001", 1047 => "11000101", 1049 => "00101111", 1050 => "10011111", 1052 => "00011011", 1053 => "11000001", 1054 => "00100111", 1055 => "10101010", 1056 => "11110011", 1057 => "11101110", 1058 => "00111011", 1060 => "01101010", 1061 => "10101100", 1062 => "00100010", 1063 => "11101000", 1065 => "11010110", 1066 => "10100001", 1067 => "00111010", 1069 => "10001110", 1071 => "01000111", 1072 => "11101101", 1074 => "11101000", 1075 => "01000110", 1077 => "00010010", 1078 => "01011011", 1079 => "10111100", 1080 => "00011001", 1081 => "00001010", 1082 => "11101010", 1084 => "01000001", 1085 => "01010001", 1087 => "01011111", 1088 => "10101101", 1092 => "11111101", 1094 => "10101000", 1095 => "00110100", 1097 => "00100100", 1098 => "10111010", 1099 => "11110001", 1100 => "11100010", 1101 => "10011111", 1102 => "11011011", 1104 => "10110010", 1105 => "01010101", 1108 => "11000110", 1109 => "10011100", 1111 => "00111110", 1112 => "00001011", 1113 => "11100000", 1115 => "00111111", 1116 => "11011000", 1118 => "01111111", 1119 => "11100011", 1121 => "01101001", 1122 => "00011101", 1123 => "11001010", 1127 => "01110101", 1128 => "00010011", 1130 => "10111010", 1133 => "00000111", 1135 => "00101000", 1136 => "10001110", 1138 => "01110001", 1141 => "11100111", 1143 => "00001010", 1144 => "01010010", 1146 => "01100000", 1147 => "01001100", 1148 => "11101010", 1149 => "10111101", 1151 => "00100111", 1152 => "01111000", 1153 => "00000001", 1157 => "11010111", 1158 => "00110101", 1159 => "10111100", 1162 => "01011000", 1164 => "11101110", 1165 => "00111111", 1166 => "10010011", 1167 => "00001110", 1169 => "01110111", 1171 => "00110101", 1173 => "10011111", 1178 => "01101010", 1179 => "11101001", 1180 => "00011111", 1181 => "00100101", 1182 => "01110000", 1183 => "10010000", 1184 => "10101000", 1185 => "11111101", 1186 => "01111000", 1187 => "10110110", 1188 => "10100010", 1189 => "01001111", 1190 => "11100101", 1191 => "11001101", 1192 => "10010010", 1193 => "10100010", 1194 => "00011011", 1198 => "10010110", 1199 => "11101101", 1200 => "10010100", 1201 => "11000011", 1202 => "00111110", 1203 => "10001010", 1205 => "10111111", 1206 => "01101111", 1207 => "00111100", 1208 => "11101011", 1209 => "10101001", 1210 => "00000100", 1211 => "11110010", 1213 => "11010011", 1214 => "10011111", 1216 => "01001101", 1218 => "11001110", 1219 => "01111000", 1220 => "00000001", 1221 => "11011011", 1223 => "11001100", 1224 => "01011011", 1226 => "00101001", 1228 => "01111010", 1229 => "10001010", 1230 => "10011011", 1232 => "00110001", 1233 => "00111000", 1235 => "11101010", 1236 => "11011111", 1237 => "11010111", 1238 => "10010000", 1239 => "10011111", 1240 => "00111111", 1241 => "10001011", 1242 => "11100010", 1243 => "11010111", 1247 => "10000001", 1248 => "11001000", 1249 => "01000111", 1250 => "00100101", 1252 => "01101001", 1253 => "00001101", 1254 => "10110110", 1255 => "10010111", 1256 => "00101101", 1257 => "01001000", 1260 => "11111001", 1261 => "01001010", 1262 => "00110110", 1263 => "11010011", 1264 => "01011111", 1265 => "00011100", 1266 => "10001010", 1267 => "11010100", 1269 => "00011000", 1270 => "10010001", 1271 => "01111010", 1272 => "10101101", 1273 => "00001100", 1275 => "10110010", 1276 => "11100010", 1278 => "11011001", 1279 => "01010111", 1280 => "01010101", 1281 => "10100010", 1282 => "01001011", 1283 => "10111010", 1285 => "10000001", 1286 => "00101100", 1287 => "00010010", 1289 => "00100001", 1290 => "00101111", 1291 => "01001011", 1292 => "01010101", 1293 => "01111100", 1294 => "00011111", 1296 => "01001101", 1297 => "11010110", 1298 => "10100110", 1299 => "11111111", 1301 => "01010101", 1302 => "11001100", 1303 => "11000000", 1305 => "00100101", 1306 => "11011000", 1307 => "11100000", 1309 => "01110000", 1310 => "00000101", 1311 => "01100010", 1312 => "00001110", 1313 => "00001000", 1314 => "01111010", 1316 => "00000101", 1317 => "11001000", 1318 => "01001100", 1320 => "00010010", 1322 => "10001100", 1324 => "10101001", 1325 => "10011110", 1328 => "00011101", 1330 => "01100000", 1331 => "10101000", 1332 => "10111001", 1335 => "01100011", 1336 => "10111101", 1337 => "10000001", 1338 => "11110111", 1339 => "01010101", 1341 => "00111111", 1342 => "11100001", 1344 => "01101110", 1345 => "00001101", 1346 => "01101011", 1347 => "11100010", 1348 => "00100010", 1349 => "01110000", 1351 => "11111101", 1352 => "11111000", 1353 => "11111110", 1355 => "11110100", 1356 => "10010110", 1359 => "11111000", 1362 => "11000011", 1363 => "10000010", 1366 => "01001100", 1367 => "01000011", 1368 => "00101011", 1369 => "11001101", 1370 => "00110110", 1371 => "10111010", 1373 => "10011010", 1374 => "11010111", 1375 => "01100011", 1377 => "10011101", 1378 => "11111110", 1379 => "10111011", 1380 => "10110100", 1381 => "00100011", 1382 => "00010010", 1383 => "01110111", 1384 => "00111100", 1385 => "11110001", 1386 => "00101101", 1387 => "10111001", 1392 => "11000110", 1393 => "10111110", 1394 => "00011111", 1395 => "00100101", 1396 => "11000000", 1399 => "11111000", 1401 => "00101101", 1402 => "00100000", 1403 => "01100001", 1404 => "00111111", 1405 => "01010011", 1407 => "01111110", 1408 => "10011001", 1410 => "01101010", 1411 => "10101010", 1412 => "00010100", 1413 => "00001110", 1414 => "10000000", 1415 => "01001110", 1416 => "00100001", 1417 => "00101101", 1418 => "11111110", 1420 => "11111101", 1421 => "00101101", 1423 => "00101001", 1424 => "00101000", 1426 => "11110100", 1427 => "10000000", 1429 => "11101010", 1430 => "01010011", 1431 => "10100010", 1433 => "11111011", 1434 => "01101100", 1435 => "11000110", 1436 => "10100100", 1437 => "00101101", 1439 => "11011110", 1440 => "10111011", 1441 => "10001001", 1443 => "00111000", 1444 => "11011100", 1449 => "10101101", 1450 => "00010100", 1452 => "11001000", 1454 => "11010000", 1455 => "01110101", 1456 => "01001000", 1457 => "00110110", 1458 => "01111110", 1459 => "11101110", 1460 => "00011000", 1464 => "00001000", 1465 => "01110101", 1466 => "11111111", 1467 => "11000101", 1469 => "11011100", 1470 => "11110011", 1473 => "00111000", 1475 => "00011001", 1477 => "00010000", 1478 => "10111001", 1479 => "01100000", 1480 => "00011011", 1481 => "00001001", 1482 => "10000001", 1483 => "00011001", 1484 => "10000010", 1485 => "01111100", 1486 => "11011011", 1488 => "00001101", 1490 => "11011011", 1491 => "00011111", 1492 => "11100011", 1493 => "00000010", 1494 => "11011100", 1495 => "01011000", 1496 => "00010101", 1497 => "01001111", 1498 => "10101001", 1499 => "01111100", 1501 => "01111001", 1503 => "11111111", 1506 => "00011100", 1507 => "01111010", 1508 => "11000100", 1509 => "10111100", 1510 => "11110111", 1511 => "11001111", 1512 => "00110011", 1514 => "10110101", 1515 => "11101111", 1516 => "01110110", 1517 => "00001000", 1518 => "00100111", 1519 => "11000100", 1520 => "11010000", 1521 => "11101011", 1524 => "10101101", 1526 => "01101100", 1527 => "00001100", 1528 => "10101100", 1529 => "00011110", 1531 => "00000110", 1532 => "11010010", 1533 => "10001001", 1534 => "01010100", 1535 => "00011111", 1537 => "01011000", 1539 => "10000001", 1540 => "10011110", 1543 => "00111101", 1544 => "00101011", 1545 => "10111110", 1547 => "00001011", 1548 => "10011110", 1551 => "11110100", 1552 => "01001011", 1553 => "01110110", 1555 => "01110110", 1556 => "00111101", 1557 => "11001100", 1559 => "10000001", 1560 => "10011000", 1561 => "11101111", 1564 => "11010101", 1566 => "01001101", 1567 => "10111101", 1568 => "00100000", 1569 => "00000110", 1571 => "10011111", 1572 => "00011110", 1573 => "01101111", 1576 => "11110001", 1577 => "01101011", 1578 => "01101100", 1579 => "01000000", 1580 => "00111001", 1581 => "01101111", 1582 => "11110000", 1583 => "01101101", 1585 => "10110000", 1587 => "00011101", 1588 => "01110001", 1589 => "10101110", 1590 => "11011100", 1592 => "11011100", 1593 => "00010110", 1594 => "11010110", 1595 => "00011110", 1596 => "11001110", 1597 => "00010100", 1598 => "00110001", 1599 => "00000110", 1600 => "10100001", 1601 => "00011110", 1602 => "01001000", 1603 => "01010100", 1604 => "10001101", 1605 => "11110000", 1606 => "01011110", 1607 => "11011001", 1608 => "10110100", 1609 => "01011111", 1610 => "00010101", 1611 => "01100011", 1613 => "01011110", 1614 => "11010110", 1615 => "01100101", 1616 => "01101111", 1617 => "10001100", 1618 => "00100101", 1619 => "11001001", 1620 => "01110101", 1621 => "11010111", 1622 => "01010000", 1623 => "01111110", 1624 => "11111001", 1625 => "10000101", 1626 => "00001110", 1627 => "00011000", 1628 => "10011010", 1630 => "01000101", 1631 => "11010000", 1632 => "01101000", 1633 => "10010011", 1634 => "01100100", 1635 => "10011001", 1636 => "00100100", 1637 => "10110011", 1638 => "00110111", 1639 => "11111011", 1640 => "10111001", 1641 => "11011100", 1642 => "00001010", 1643 => "10101010", 1645 => "10010011", 1648 => "01100000", 1649 => "01111111", 1652 => "11111101", 1653 => "11010110", 1654 => "00100101", 1655 => "11000100", 1657 => "10101110", 1658 => "11101110", 1659 => "00101100", 1660 => "01000001", 1662 => "00110110", 1663 => "11010011", 1664 => "11000011", 1665 => "10011111", 1666 => "10011001", 1667 => "01000001", 1668 => "10101010", 1669 => "01100110", 1670 => "10011000", 1671 => "00100001", 1672 => "10101011", 1678 => "00000100", 1680 => "11100011", 1681 => "01101100", 1682 => "01001110", 1683 => "11111100", 1686 => "01010111", 1687 => "10100010", 1689 => "00111001", 1690 => "00001101", 1692 => "11000000", 1693 => "01100100", 1694 => "01010001", 1696 => "10010000", 1697 => "01010111", 1698 => "11100011", 1699 => "11101101", 1700 => "11111101", 1701 => "11000011", 1702 => "01111011", 1703 => "11001110", 1704 => "11111011", 1706 => "00101000", 1707 => "11001111", 1708 => "01111110", 1709 => "00000011", 1710 => "00101011", 1711 => "00101111", 1712 => "10000010", 1713 => "01100101", 1715 => "00111001", 1716 => "10111101", 1717 => "11101011", 1718 => "10101000", 1719 => "00011110", 1721 => "01111111", 1722 => "10001010", 1723 => "11000101", 1724 => "11111110", 1726 => "01001010", 1727 => "01010001", 1729 => "10011000", 1730 => "00111000", 1731 => "00110111", 1732 => "00001110", 1735 => "01101001", 1737 => "10101111", 1738 => "01000010", 1739 => "01000101", 1740 => "01110000", 1742 => "11100010", 1743 => "01000011", 1744 => "11000101", 1745 => "00100111", 1746 => "01010101", 1748 => "01011101", 1749 => "01001000", 1752 => "10111011", 1753 => "11011111", 1754 => "00011001", 1756 => "00000001", 1758 => "00101010", 1759 => "00000010", 1760 => "01001101", 1761 => "10011111", 1763 => "10010011", 1764 => "10111011", 1765 => "00110110", 1766 => "11101010", 1767 => "01101100", 1769 => "10000010", 1770 => "00011011", 1771 => "00110111", 1772 => "01100101", 1773 => "10101010", 1775 => "11101100", 1777 => "11100001", 1778 => "00111110", 1779 => "01000010", 1780 => "11010000", 1781 => "00110110", 1782 => "00101010", 1783 => "01110000", 1784 => "00111111", 1785 => "00101110", 1786 => "11011110", 1788 => "10110110", 1789 => "10001111", 1790 => "10011001", 1792 => "10001000", 1793 => "01001011", 1795 => "01010100", 1796 => "01100101", 1797 => "11011011", 1798 => "10110010", 1799 => "01010000", 1800 => "11011010", 1801 => "00001101", 1802 => "10001001", 1803 => "00011010", 1805 => "11011000", 1809 => "00100011", 1810 => "11101110", 1811 => "10110110", 1812 => "00101111", 1813 => "10111101", 1814 => "11001111", 1815 => "10010000", 1817 => "11100001", 1818 => "10010111", 1819 => "11100001", 1820 => "10101100", 1821 => "10001111", 1824 => "11110000", 1825 => "00001001", 1826 => "10111011", 1827 => "01111000", 1828 => "10011111", 1829 => "11000110", 1832 => "01001100", 1833 => "01000100", 1835 => "01000100", 1836 => "11111100", 1837 => "10101011", 1840 => "11111110", 1841 => "11110000", 1842 => "01000001", 1843 => "00101011", 1844 => "10001001", 1845 => "11100010", 1846 => "11000001", 1847 => "00000001", 1848 => "10111100", 1849 => "00000110", 1850 => "00110001", 1853 => "10011010", 1854 => "01010011", 1855 => "00110000", 1856 => "11000101", 1857 => "11100101", 1858 => "11111010", 1859 => "00010001", 1860 => "11110010", 1862 => "01011011", 1863 => "10101111", 1864 => "10000101", 1866 => "00111111", 1868 => "11101011", 1871 => "10111101", 1872 => "00010001", 1873 => "10001100", 1874 => "11000001", 1875 => "01100001", 1876 => "00000001", 1877 => "11001100", 1878 => "00110001", 1879 => "00110010", 1882 => "01110101", 1883 => "10011110", 1884 => "10010110", 1885 => "00100100", 1887 => "11101100", 1888 => "11010100", 1890 => "10111001", 1891 => "10011011", 1893 => "11111000", 1894 => "10111001", 1895 => "01100001", 1896 => "10111110", 1897 => "11001100", 1899 => "00000111", 1901 => "11111011", 1902 => "11111000", 1903 => "10011110", 1904 => "11010010", 1905 => "00110110", 1906 => "00010001", 1907 => "10110110", 1908 => "10001001", 1909 => "10001101", 1910 => "00000010", 1911 => "11000011", 1912 => "11001111", 1914 => "11110100", 1916 => "00100010", 1917 => "10001110", 1919 => "11111111", 1920 => "00110010", 1921 => "00101001", 1927 => "10001001", 1928 => "10101010", 1930 => "10001010", 1932 => "01100111", 1933 => "11001111", 1934 => "01010011", 1935 => "11101000", 1937 => "01110110", 1938 => "00001101", 1939 => "11110101", 1940 => "00111111", 1941 => "01110001", 1942 => "10101100", 1945 => "11101000", 1946 => "11000011", 1947 => "11100101", 1948 => "11111100", 1949 => "10101011", 1951 => "01010100", 1952 => "10010011", 1954 => "11100100", 1955 => "00000111", 1958 => "00011110", 1959 => "00010001", 1960 => "11111111", 1961 => "10011100", 1962 => "01101000", 1966 => "11111010", 1967 => "01001000", 1968 => "11111101", 1970 => "01110001", 1971 => "10110010", 1973 => "00110101", 1975 => "10001100", 1976 => "01010000", 1977 => "01010011", 1980 => "01001001", 1981 => "10101000", 1982 => "00011011", 1983 => "11010011", 1984 => "10101110", 1985 => "01111101", 1988 => "01011100", 1989 => "01000101", 1992 => "11111111", 1993 => "01000011", 1994 => "11010100", 1998 => "11111100", 2000 => "11010010", 2001 => "01000110", 2002 => "00101101", 2003 => "01011001", 2006 => "00001010", 2007 => "10000001", 2009 => "10110000", 2010 => "01111100", 2011 => "10000110", 2012 => "01111001", 2014 => "00100111", 2015 => "01111001", 2016 => "11001010", 2017 => "00011011", 2018 => "00110001", 2019 => "00000100", 2020 => "10000000", 2021 => "00101010", 2022 => "10101111", 2023 => "00111101", 2024 => "11100111", 2025 => "00000111", 2027 => "00011011", 2028 => "11000001", 2030 => "00000010", 2031 => "10110110", 2032 => "11001000", 2034 => "10111111", 2035 => "01101011", 2037 => "00010010", 2038 => "10000011", 2039 => "10010111", 2040 => "11100101", 2041 => "01010000", 2044 => "01111001", 2046 => "11100010", 2047 => "11100100", 2049 => "00011111", 2051 => "01101101", 2052 => "00000101", 2053 => "00110101", 2054 => "00000100", 2056 => "00001000", 2057 => "00111010", 2059 => "10110101", 2060 => "11010110", 2061 => "01000100", 2062 => "00100000", 2064 => "01111110", 2065 => "11110000", 2066 => "11110001", 2067 => "11000000", 2068 => "10110101", 2070 => "11110000", 2071 => "11100110", 2072 => "01110010", 2075 => "11010111", 2076 => "10010001", 2077 => "10010010", 2078 => "00101101", 2079 => "00110110", 2081 => "00001000", 2082 => "00011000", 2083 => "01010000", 2085 => "01110010", 2086 => "00001001", 2091 => "10001001", 2093 => "10111010", 2094 => "00011110", 2095 => "11001010", 2096 => "10010110", 2098 => "10101100", 2099 => "01110101", 2101 => "11110101", 2102 => "10100100", 2103 => "00011000", 2104 => "00100010", 2106 => "11101110", 2107 => "10001111", 2108 => "11111010", 2109 => "10001100", 2110 => "11111011", 2111 => "11110010", 2112 => "01001101", 2114 => "11111000", 2116 => "00100111", 2117 => "01100100", 2118 => "01001101", 2119 => "11001000", 2120 => "11110010", 2121 => "01111110", 2122 => "01010101", 2123 => "00010000", 2125 => "00101100", 2126 => "00010111", 2128 => "01001001", 2130 => "01101111", 2132 => "10110011", 2133 => "10110001", 2136 => "11001010", 2137 => "00010110", 2138 => "00111000", 2139 => "00011000", 2140 => "10010111", 2142 => "00111101", 2144 => "01110100", 2146 => "01010111", 2147 => "10101010", 2149 => "10100101", 2151 => "10001100", 2152 => "11110100", 2153 => "01000001", 2154 => "01000000", 2155 => "00001000", 2158 => "10100111", 2160 => "11100101", 2161 => "00100111", 2162 => "00111010", 2163 => "11101110", 2166 => "01011110", 2167 => "10000110", 2168 => "10111100", 2169 => "00001001", 2171 => "00101101", 2172 => "11000101", 2174 => "11100100", 2175 => "01001111", 2177 => "01101010", 2178 => "01110100", 2179 => "10001001", 2180 => "00010110", 2182 => "10110100", 2183 => "01010111", 2184 => "10011100", 2186 => "00011010", 2187 => "10111000", 2188 => "10111100", 2191 => "10000111", 2193 => "01001011", 2194 => "00111110", 2196 => "00100011", 2197 => "11011111", 2199 => "10110101", 2200 => "01111011", 2202 => "11111000", 2204 => "01101100", 2206 => "00010110", 2207 => "10111000", 2208 => "11011010", 2209 => "11111100", 2210 => "11100111", 2211 => "01101000", 2212 => "11100011", 2213 => "11111110", 2214 => "11101011", 2216 => "10001100", 2218 => "10110001", 2219 => "10110011", 2221 => "10000110", 2224 => "11110001", 2225 => "00000010", 2226 => "00000110", 2227 => "10001011", 2228 => "10100010", 2229 => "01110110", 2230 => "00000110", 2233 => "11000100", 2234 => "11101111", 2235 => "11011100", 2236 => "00001111", 2237 => "00010110", 2238 => "00011000", 2239 => "00111010", 2240 => "01111010", 2242 => "01111111", 2243 => "00101111", 2244 => "10111101", 2246 => "01111101", 2247 => "11010101", 2248 => "11001100", 2250 => "01011111", 2251 => "10011000", 2252 => "10010111", 2253 => "01010010", 2255 => "10010110", 2256 => "10101001", 2257 => "10011001", 2258 => "00011001", 2261 => "10111111", 2262 => "10111000", 2264 => "00001110", 2265 => "01000111", 2267 => "01111110", 2268 => "10010000", 2269 => "00101111", 2270 => "11111001", 2271 => "10110100", 2272 => "00111011", 2273 => "10101111", 2275 => "00101110", 2276 => "00011011", 2277 => "01000010", 2279 => "10100010", 2280 => "00010010", 2281 => "10110100", 2282 => "10111101", 2285 => "11111101", 2286 => "10100010", 2287 => "01011001", 2289 => "01010011", 2291 => "10101110", 2293 => "01111000", 2296 => "01011111", 2298 => "00000100", 2299 => "00000101", 2300 => "01111010", 2301 => "11011001", 2302 => "01001101", 2303 => "00101111", 2304 => "00111010", 2305 => "10110110", 2306 => "11001011", 2309 => "00010011", 2311 => "10001101", 2312 => "10000011", 2313 => "01001110", 2315 => "10010100", 2317 => "10100101", 2320 => "10111000", 2321 => "10100010", 2324 => "11110010", 2325 => "01000010", 2326 => "00000101", 2328 => "11110010", 2329 => "01000100", 2330 => "11010011", 2331 => "01111011", 2333 => "01101110", 2334 => "01010110", 2336 => "00000001", 2337 => "01011000", 2338 => "01100111", 2340 => "01110100", 2341 => "11100101", 2343 => "11101001", 2345 => "11111101", 2346 => "10011101", 2347 => "00111000", 2349 => "00110111", 2352 => "01010110", 2354 => "01101011", 2355 => "11011001", 2356 => "00010100", 2357 => "00101010", 2359 => "00111110", 2360 => "10110001", 2361 => "01101000", 2363 => "00011110", 2364 => "10001101", 2365 => "01001011", 2366 => "00011000", 2367 => "01101110", 2368 => "11001010", 2369 => "10001100", 2371 => "11101110", 2374 => "01110110", 2376 => "00100101", 2378 => "11111010", 2379 => "11111000", 2380 => "11000111", 2381 => "11000110", 2383 => "01010111", 2384 => "11101011", 2385 => "01101100", 2386 => "00100111", 2387 => "01111101", 2389 => "00011101", 2391 => "00101110", 2392 => "10110000", 2393 => "10010100", 2394 => "11100010", 2395 => "01001011", 2396 => "00001010", 2397 => "10011000", 2398 => "01100100", 2400 => "00010010", 2403 => "10001101", 2405 => "11001100", 2407 => "11101100", 2408 => "00000001", 2410 => "10001011", 2411 => "10010101", 2412 => "11110001", 2413 => "01010101", 2414 => "10111110", 2415 => "11111101", 2416 => "11011000", 2417 => "10100101", 2418 => "11010010", 2419 => "11100000", 2420 => "00100101", 2421 => "10101011", 2422 => "00101011", 2423 => "01011010", 2425 => "10001100", 2427 => "11001111", 2428 => "10001110", 2431 => "01110101", 2434 => "00010111", 2436 => "00010110", 2437 => "11010111", 2438 => "11111111", 2439 => "11010110", 2440 => "00111100", 2445 => "11101110", 2447 => "01001000", 2448 => "11111111", 2449 => "11010001", 2450 => "01010101", 2452 => "11001001", 2453 => "01100101", 2455 => "01100011", 2456 => "00011100", 2457 => "11001010", 2458 => "11100010", 2459 => "01101111", 2460 => "11111111", 2461 => "01010100", 2462 => "10011110", 2463 => "10011101", 2464 => "01111110", 2465 => "01110001", 2466 => "10010000", 2467 => "01000100", 2468 => "00001001", 2469 => "10100001", 2470 => "00011111", 2471 => "01110011", 2472 => "11100011", 2473 => "11110010", 2474 => "11000110", 2475 => "11101011", 2476 => "10000100", 2477 => "00001001", 2478 => "10100000", 2479 => "11011010", 2480 => "00000011", 2481 => "10111100", 2482 => "01001011", 2483 => "10010010", 2484 => "11101001", 2485 => "10000101", 2489 => "00001100", 2491 => "00110111", 2492 => "01111000", 2493 => "00110100", 2494 => "10100111", 2495 => "10110100", 2497 => "00110110", 2498 => "10111010", 2499 => "11111000", 2500 => "00100100", 2501 => "01001000", 2503 => "11111110", 2504 => "10110010", 2505 => "10010000", 2506 => "11011010", 2507 => "00111001", 2508 => "10100110", 2509 => "00010001", 2511 => "11010011", 2512 => "00110010", 2513 => "01111110", 2514 => "01011001", 2516 => "11100001", 2517 => "00101111", 2520 => "01100010", 2526 => "11000001", 2528 => "10111110", 2530 => "01101001", 2531 => "11110011", 2532 => "10011011", 2533 => "01010111", 2534 => "11000011", 2535 => "11111011", 2537 => "01100011", 2538 => "01101010", 2540 => "10100000", 2541 => "10010101", 2542 => "11100001", 2543 => "00001000", 2544 => "10101100", 2546 => "01101111", 2547 => "11011100", 2548 => "01100100", 2549 => "00001111", 2550 => "00000011", 2551 => "01000111", 2553 => "10000101", 2555 => "10100011", 2556 => "10001000", 2558 => "10000000", 2559 => "10100110", 2562 => "00101101", 2563 => "00010110", 2564 => "01110010", 2565 => "01110001", 2566 => "11111011", 2567 => "00100010", 2568 => "00111111", 2570 => "10011001", 2571 => "00100001", 2573 => "01011001", 2574 => "00010101", 2575 => "00100101", 2578 => "01001011", 2579 => "01111011", 2580 => "00000001", 2581 => "01101001", 2582 => "00110101", 2583 => "00011000", 2584 => "00011101", 2586 => "00100000", 2589 => "11010011", 2590 => "00111101", 2591 => "00001011", 2594 => "10101101", 2595 => "10010101", 2596 => "00000111", 2597 => "01100100", 2598 => "10000001", 2599 => "10110011", 2600 => "11001001", 2601 => "10111010", 2602 => "01000010", 2603 => "11111111", 2604 => "01011100", 2606 => "01001010", 2607 => "10000111", 2608 => "11001010", 2609 => "01001001", 2611 => "01100010", 2612 => "11110000", 2613 => "00011100", 2614 => "00001010", 2615 => "00001010", 2617 => "11000110", 2618 => "10011111", 2619 => "11101001", 2620 => "01011001", 2622 => "01110010", 2623 => "01100011", 2624 => "01110001", 2625 => "00011111", 2626 => "00101101", 2629 => "01000100", 2630 => "11101100", 2631 => "00011100", 2632 => "00011011", 2635 => "00110011", 2636 => "01011011", 2637 => "10000111", 2640 => "00111000", 2641 => "10111111", 2643 => "10110100", 2644 => "00101000", 2646 => "11001010", 2648 => "11000101", 2650 => "00100100", 2651 => "11100010", 2652 => "01100011", 2653 => "11000110", 2654 => "00110100", 2655 => "10110110", 2656 => "10011100", 2657 => "11100010", 2658 => "01011011", 2659 => "10010000", 2660 => "00000100", 2661 => "10111110", 2662 => "00000001", 2664 => "11100011", 2665 => "10110000", 2666 => "10100001", 2667 => "11001011", 2668 => "11110011", 2671 => "01011010", 2672 => "00001001", 2673 => "01001111", 2674 => "11010110", 2675 => "10010011", 2676 => "11101001", 2679 => "01111010", 2681 => "00000011", 2682 => "01001101", 2683 => "10011110", 2685 => "00100001", 2686 => "11010100", 2687 => "00011111", 2688 => "01000011", 2690 => "01000011", 2691 => "11100001", 2692 => "11100011", 2693 => "10101111", 2695 => "10101101", 2697 => "10110011", 2698 => "11011011", 2699 => "01010010", 2700 => "01001011", 2701 => "10100011", 2702 => "11010100", 2704 => "10111010", 2705 => "00110011", 2707 => "00001101", 2708 => "11111101", 2709 => "11100000", 2710 => "10010001", 2711 => "00010001", 2712 => "10001010", 2714 => "11010101", 2715 => "11111001", 2717 => "11100100", 2718 => "01111010", 2719 => "11001001", 2720 => "01110000", 2721 => "00010100", 2722 => "11011111", 2723 => "01000000", 2724 => "10101111", 2726 => "01100100", 2728 => "00111111", 2729 => "00111000", 2731 => "01011101", 2732 => "00001101", 2733 => "10111010", 2736 => "01111001", 2737 => "10010110", 2740 => "00110111", 2744 => "11101000", 2749 => "10010100", 2750 => "01110010", 2752 => "01100111", 2755 => "11011000", 2757 => "11010010", 2758 => "10011001", 2759 => "10001111", 2761 => "00010100", 2762 => "10100010", 2764 => "00000110", 2766 => "11010011", 2767 => "10001101", 2768 => "10001000", 2771 => "11001000", 2772 => "00010001", 2773 => "10101111", 2774 => "01010011", 2776 => "11011000", 2778 => "11101111", 2779 => "11010111", 2780 => "11101101", 2781 => "10011001", 2782 => "10010111", 2783 => "11100110", 2784 => "11100110", 2785 => "01101101", 2786 => "10101110", 2787 => "10010011", 2789 => "11101011", 2790 => "01011011", 2791 => "11011110", 2792 => "00011111", 2793 => "00001010", 2794 => "10011100", 2795 => "00000001", 2796 => "10110110", 2798 => "11110111", 2799 => "00110011", 2802 => "00110000", 2803 => "10100100", 2808 => "10000110", 2809 => "01010100", 2810 => "10111100", 2814 => "01100100", 2815 => "00100101", 2816 => "10101010", 2817 => "00000101", 2818 => "10111110", 2819 => "10001000", 2821 => "01110111", 2824 => "11100000", 2827 => "10101010", 2829 => "11100111", 2831 => "01010001", 2832 => "10011011", 2833 => "00010110", 2836 => "11011111", 2837 => "00110101", 2838 => "00000100", 2839 => "10010011", 2840 => "10000111", 2842 => "10001110", 2843 => "00001011", 2845 => "11100111", 2846 => "11110001", 2847 => "10101110", 2848 => "11011111", 2849 => "00111001", 2851 => "00101111", 2852 => "11101000", 2853 => "11001000", 2855 => "11010001", 2856 => "00110110", 2857 => "11011101", 2858 => "00100100", 2859 => "01000001", 2861 => "11111101", 2862 => "11001000", 2863 => "11011110", 2866 => "11000011", 2867 => "11100011", 2869 => "11011011", 2870 => "11011000", 2871 => "11001100", 2872 => "10101010", 2874 => "00000110", 2875 => "01100010", 2878 => "00000111", 2879 => "01101100", 2880 => "01001000", 2881 => "11010010", 2882 => "11111011", 2883 => "00110000", 2885 => "01000011", 2886 => "10011100", 2888 => "10100000", 2889 => "11101110", 2890 => "00011000", 2892 => "01110111", 2895 => "10010001", 2896 => "01100111", 2898 => "00110111", 2900 => "01000101", 2901 => "10101001", 2903 => "10111110", 2906 => "00000010", 2907 => "11010101", 2908 => "01111011", 2909 => "00011100", 2910 => "01101111", 2911 => "11011000", 2912 => "00001100", 2916 => "10000100", 2917 => "11110110", 2918 => "00011001", 2919 => "00001100", 2920 => "00100100", 2921 => "01011011", 2922 => "10110001", 2923 => "01111011", 2924 => "10101110", 2925 => "00001010", 2926 => "10011011", 2927 => "00101100", 2928 => "01001100", 2929 => "11111100", 2930 => "00110110", 2931 => "11010100", 2932 => "10110110", 2933 => "00001101", 2935 => "11110101", 2936 => "10101110", 2938 => "10101000", 2939 => "01010000", 2940 => "11001010", 2941 => "01001100", 2943 => "01111110", 2945 => "01010110", 2946 => "01110111", 2947 => "00111011", 2948 => "11000011", 2949 => "11110100", 2951 => "00010110", 2952 => "00001000", 2953 => "10011101", 2954 => "01100011", 2955 => "01100001", 2956 => "10000000", 2958 => "10110110", 2959 => "01101111", 2961 => "11011110", 2962 => "11111111", 2963 => "10111010", 2964 => "01010100", 2966 => "10001011", 2967 => "10101000", 2970 => "11111100", 2972 => "11010011", 2973 => "11100010", 2975 => "00001110", 2976 => "00000001", 2977 => "10110100", 2978 => "10111000", 2980 => "00100001", 2983 => "10011110", 2984 => "00011100", 2985 => "00110101", 2986 => "00000100", 2988 => "11100000", 2989 => "01111011", 2990 => "11011000", 2992 => "11101000", 2993 => "00101110", 2994 => "11101100", 2995 => "10001001", 2997 => "00111001", 2999 => "11011011", 3001 => "01111101", 3002 => "11000011", 3004 => "01110111", 3005 => "01000010", 3006 => "01101101", 3008 => "00101000", 3011 => "11001000", 3014 => "01010011", 3016 => "00111010", 3018 => "00010010", 3021 => "01010000", 3022 => "11100110", 3023 => "01001100", 3024 => "10011000", 3028 => "01111100", 3031 => "11000001", 3032 => "10001111", 3033 => "01010101", 3034 => "00101000", 3038 => "10000101", 3039 => "00001001", 3040 => "00011110", 3041 => "10011111", 3045 => "01001101", 3048 => "01010100", 3049 => "10010100", 3050 => "10101101", 3053 => "01100010", 3054 => "01111010", 3055 => "01101101", 3057 => "11100111", 3058 => "01010001", 3061 => "11100110", 3062 => "01000111", 3063 => "10110011", 3064 => "10100000", 3065 => "01000011", 3066 => "11100011", 3067 => "10110001", 3068 => "00101001", 3069 => "11101001", 3070 => "11110111", 3071 => "00011111", 3072 => "01001110", 3073 => "00110101", 3079 => "11110110", 3080 => "11000010", 3081 => "11010000", 3082 => "00101100", 3083 => "01100101", 3084 => "11101010", 3085 => "11011000", 3089 => "01111010", 3090 => "11000010", 3091 => "00101001", 3092 => "11011111", 3094 => "11000000", 3095 => "11110100", 3096 => "11101111", 3098 => "01011010", 3100 => "10000000", 3102 => "01000111", 3103 => "10001100", 3104 => "01101101", 3105 => "11111110", 3106 => "10010011", 3107 => "01111101", 3109 => "10001101", 3110 => "01100101", 3111 => "11100100", 3112 => "11100011", 3113 => "11100110", 3115 => "01011111", 3116 => "10110000", 3117 => "00111010", 3119 => "11000110", 3120 => "10011110", 3121 => "11001110", 3122 => "10011011", 3123 => "01110111", 3124 => "11010100", 3125 => "01011001", 3129 => "00101001", 3131 => "11011101", 3132 => "00110000", 3133 => "01110000", 3134 => "00111001", 3135 => "11001100", 3136 => "11001101", 3139 => "10010100", 3140 => "00110011", 3141 => "11001100", 3142 => "01001001", 3144 => "10010110", 3146 => "00111110", 3147 => "10000011", 3148 => "00110101", 3149 => "01110000", 3150 => "01011000", 3151 => "00011010", 3152 => "10001100", 3154 => "00111011", 3155 => "10111100", 3156 => "01110000", 3157 => "00110010", 3158 => "11100101", 3159 => "00111000", 3160 => "11100010", 3161 => "00111000", 3162 => "10000111", 3163 => "01001001", 3165 => "10000011", 3166 => "00101100", 3168 => "11001001", 3169 => "00100111", 3172 => "01101000", 3173 => "01110011", 3175 => "10011010", 3176 => "00110011", 3177 => "11100100", 3178 => "11101111", 3179 => "11010101", 3180 => "01011001", 3181 => "11010101", 3182 => "10110001", 3184 => "10010011", 3185 => "00110000", 3187 => "00011011", 3188 => "10100110", 3189 => "10100011", 3192 => "01110101", 3193 => "10100000", 3195 => "01001101", 3196 => "10000001", 3197 => "11010101", 3199 => "01011010", 3200 => "11010001", 3201 => "10010100", 3202 => "10111011", 3205 => "01010101", 3206 => "01110110", 3207 => "11100101", 3208 => "01011100", 3209 => "00000100", 3210 => "00101100", 3211 => "00100010", 3212 => "00000111", 3213 => "01110110", 3214 => "10111001", 3215 => "11000010", 3216 => "11111111", 3217 => "00101101", 3218 => "01111001", 3219 => "01010011", 3220 => "01110010", 3222 => "11011111", 3223 => "10110011", 3226 => "11101111", 3227 => "11100111", 3228 => "00011010", 3229 => "01001100", 3230 => "11111000", 3232 => "00110000", 3233 => "10001010", 3235 => "00110000", 3237 => "10011010", 3239 => "10111100", 3240 => "11100110", 3242 => "11011111", 3243 => "00111010", 3244 => "10111100", 3246 => "00010100", 3247 => "00000010", 3248 => "10100100", 3249 => "01011100", 3250 => "00101011", 3251 => "00000010", 3254 => "10100010", 3256 => "11101010", 3257 => "10101110", 3258 => "11111010", 3259 => "10001000", 3261 => "11010111", 3263 => "01100011", 3267 => "11010001", 3268 => "01000111", 3271 => "00100110", 3272 => "11010010", 3273 => "01000100", 3274 => "11110110", 3275 => "00101000", 3276 => "01010011", 3277 => "01010101", 3279 => "10101100", 3280 => "00110100", 3281 => "10000010", 3282 => "00111110", 3284 => "10101001", 3285 => "01011111", 3286 => "10101100", 3287 => "10010100", 3288 => "00011111", 3289 => "10011100", 3291 => "11010011", 3292 => "00001101", 3295 => "01011011", 3296 => "11000001", 3298 => "10011000", 3300 => "00110110", 3301 => "10000011", 3302 => "10110010", 3303 => "10001000", 3304 => "11010111", 3307 => "11010000", 3308 => "01101111", 3309 => "10110101", 3310 => "11011010", 3311 => "00011011", 3312 => "00110110", 3313 => "10001111", 3314 => "00001111", 3317 => "11001000", 3318 => "10000010", 3319 => "10101111", 3321 => "10001011", 3322 => "00000010", 3323 => "00001000", 3326 => "11101011", 3327 => "00011101", 3329 => "11010100", 3331 => "10111011", 3333 => "10111010", 3334 => "11111001", 3335 => "10010000", 3337 => "01010011", 3339 => "01100100", 3340 => "01111010", 3342 => "11010011", 3343 => "11110001", 3344 => "10101010", 3345 => "10010010", 3346 => "00110010", 3347 => "10101111", 3348 => "00101010", 3350 => "10100111", 3351 => "11110111", 3352 => "01010111", 3353 => "01000011", 3354 => "10010101", 3355 => "00001010", 3356 => "10000000", 3357 => "00111010", 3358 => "00000011", 3361 => "01010011", 3362 => "01111110", 3363 => "00110100", 3364 => "00011111", 3365 => "11111001", 3366 => "11101101", 3367 => "11101010", 3369 => "00010111", 3373 => "11001100", 3375 => "01010001", 3377 => "10101100", 3378 => "00110100", 3379 => "00010111", 3380 => "10111101", 3381 => "10010000", 3382 => "11011101", 3383 => "00011001", 3384 => "11010001", 3385 => "00110010", 3386 => "10110011", 3388 => "01010010", 3391 => "01100101", 3392 => "01001110", 3393 => "10000011", 3395 => "11000000", 3397 => "10111111", 3398 => "01010111", 3399 => "10010000", 3400 => "10010101", 3401 => "11010010", 3402 => "10101011", 3404 => "01010111", 3405 => "01010111", 3406 => "11101010", 3407 => "11011111", 3408 => "00100001", 3412 => "10001010", 3413 => "10011000", 3414 => "00101111", 3416 => "10111001", 3418 => "01100001", 3419 => "11010010", 3420 => "01101010", 3421 => "01010001", 3422 => "11111001", 3423 => "11101010", 3424 => "01100111", 3425 => "01010011", 3426 => "10000011", 3427 => "10100000", 3428 => "11100100", 3430 => "01010011", 3431 => "11011010", 3432 => "00111101", 3433 => "10111111", 3434 => "10110001", 3436 => "01000011", 3437 => "01000110", 3438 => "11001110", 3439 => "11010011", 3440 => "00101101", 3441 => "11111100", 3442 => "01001011", 3443 => "00001110", 3444 => "10001101", 3445 => "00001010", 3446 => "00011010", 3447 => "11100110", 3449 => "00110100", 3450 => "01000011", 3453 => "10111001", 3454 => "00011111", 3455 => "10011100", 3457 => "01011110", 3459 => "11100010", 3460 => "00011101", 3461 => "00101011", 3462 => "01100000", 3463 => "01110111", 3467 => "01100101", 3470 => "01111010", 3472 => "01100110", 3473 => "00000100", 3474 => "10101110", 3475 => "10101110", 3476 => "11100110", 3478 => "01001010", 3480 => "11110111", 3481 => "11111010", 3483 => "11110011", 3484 => "00100100", 3485 => "11010101", 3486 => "11111001", 3487 => "10101100", 3489 => "11111011", 3490 => "01011001", 3494 => "00110000", 3495 => "10010111", 3496 => "10110101", 3497 => "01111010", 3499 => "00011001", 3501 => "10111011", 3502 => "01010000", 3503 => "10000001", 3504 => "00000010", 3505 => "01010001", 3506 => "00111101", 3507 => "10011001", 3509 => "11000110", 3510 => "00001110", 3512 => "10101110", 3513 => "11011010", 3515 => "00111100", 3516 => "01100110", 3518 => "11000001", 3519 => "01011011", 3520 => "00000100", 3521 => "01110100", 3523 => "00011111", 3524 => "00111110", 3525 => "10001101", 3526 => "00100100", 3527 => "00001000", 3528 => "00110000", 3529 => "00110101", 3530 => "01110111", 3532 => "10000100", 3534 => "01100100", 3535 => "10000101", 3536 => "01000100", 3537 => "11011011", 3538 => "01000101", 3539 => "10101110", 3540 => "10010010", 3541 => "01010001", 3542 => "10010110", 3543 => "10010111", 3547 => "11000101", 3549 => "10111000", 3550 => "11111100", 3554 => "10010111", 3556 => "01111100", 3557 => "00011111", 3558 => "01001100", 3560 => "01110011", 3563 => "01110100", 3564 => "10100001", 3565 => "11010000", 3566 => "00011100", 3567 => "01111110", 3568 => "11100010", 3570 => "01000001", 3571 => "00010101", 3572 => "00001000", 3573 => "01000011", 3574 => "01010000", 3575 => "10100111", 3576 => "00100100", 3577 => "01101011", 3580 => "00011100", 3581 => "00001110", 3582 => "11000010", 3583 => "10100011", 3584 => "11100010", 3588 => "01110101", 3589 => "00100111", 3591 => "10100111", 3593 => "00011101", 3595 => "01000001", 3596 => "00001101", 3597 => "11111111", 3601 => "00000011", 3602 => "10010011", 3603 => "11100001", 3604 => "01001100", 3606 => "10010101", 3607 => "11100110", 3609 => "01110011", 3613 => "01111011", 3614 => "10000000", 3615 => "10111100", 3616 => "01010110", 3618 => "00000010", 3619 => "11001011", 3621 => "10111111", 3622 => "11000010", 3623 => "01001011", 3624 => "11000000", 3625 => "01001111", 3626 => "00110110", 3628 => "11100111", 3631 => "01110110", 3632 => "10110101", 3634 => "00110000", 3635 => "11001011", 3636 => "00110101", 3637 => "10010100", 3638 => "00001001", 3639 => "10110101", 3644 => "10101111", 3645 => "01101001", 3647 => "00111001", 3648 => "10001101", 3649 => "00111011", 3650 => "00000101", 3651 => "00101001", 3652 => "11000110", 3654 => "00010011", 3656 => "10000110", 3658 => "11100000", 3659 => "10111100", 3660 => "00101110", 3662 => "00010000", 3663 => "00111100", 3664 => "00111011", 3665 => "10111010", 3668 => "11001001", 3670 => "10011001", 3671 => "01010111", 3672 => "01010011", 3675 => "10111111", 3676 => "01000110", 3677 => "01000001", 3679 => "11000011", 3680 => "00100000", 3681 => "01101100", 3683 => "11101100", 3684 => "10011001", 3685 => "11001001", 3686 => "00011110", 3690 => "01110001", 3691 => "01011100", 3692 => "01011101", 3693 => "00010000", 3694 => "11001101", 3695 => "11111000", 3696 => "00001000", 3697 => "11010101", 3700 => "00100100", 3701 => "10110101", 3702 => "10001101", 3703 => "00011101", 3705 => "01100110", 3706 => "10110001", 3707 => "01010110", 3708 => "01110110", 3709 => "11110110", 3710 => "01110100", 3713 => "10101100", 3715 => "00100111", 3716 => "11000000", 3717 => "01010001", 3719 => "11011010", 3720 => "01000010", 3722 => "01001000", 3724 => "01000010", 3726 => "11011101", 3727 => "01101010", 3729 => "11111100", 3732 => "00111001", 3734 => "10011110", 3735 => "01000011", 3736 => "01111110", 3737 => "00010111", 3739 => "00011000", 3740 => "11111110", 3743 => "11010110", 3746 => "10100100", 3749 => "00010110", 3752 => "01101010", 3753 => "11111010", 3755 => "01111010", 3756 => "01010011", 3757 => "10010101", 3758 => "00111100", 3759 => "01101011", 3761 => "11010011", 3762 => "01001111", 3763 => "00010011", 3764 => "11011101", 3767 => "11100110", 3768 => "10011000", 3770 => "01000111", 3771 => "00001000", 3772 => "01000000", 3773 => "01101111", 3774 => "01000010", 3775 => "10101110", 3777 => "10110001", 3778 => "00000110", 3781 => "01101010", 3784 => "11011111", 3785 => "00110101", 3786 => "00101101", 3787 => "10111111", 3788 => "11000000", 3790 => "00111000", 3792 => "00100100", 3793 => "11001010", 3794 => "01000010", 3795 => "10111000", 3796 => "11101000", 3797 => "01101111", 3798 => "01001000", 3800 => "10001001", 3801 => "10111001", 3802 => "10000010", 3803 => "10100011", 3804 => "10111100", 3805 => "01110101", 3806 => "00100010", 3807 => "10111011", 3808 => "01110100", 3809 => "11001010", 3811 => "11010000", 3812 => "11100100", 3813 => "00001110", 3814 => "10010101", 3815 => "01111001", 3816 => "01111011", 3817 => "01011010", 3818 => "11010001", 3819 => "00110111", 3820 => "11111001", 3821 => "10000000", 3822 => "00100001", 3823 => "10100111", 3824 => "01110111", 3825 => "11111011", 3826 => "10111100", 3828 => "11100100", 3829 => "00111100", 3830 => "01101101", 3832 => "11110000", 3833 => "01101101", 3834 => "10111111", 3835 => "00001001", 3836 => "01000111", 3837 => "10011010", 3840 => "11101000", 3841 => "11001101", 3843 => "11000001", 3844 => "11010100", 3846 => "00101010", 3849 => "11001110", 3850 => "00110111", 3851 => "01001011", 3852 => "01011010", 3853 => "01000001", 3854 => "10010101", 3855 => "11100000", 3856 => "10100011", 3860 => "11010001", 3862 => "00110101", 3863 => "11011001", 3865 => "00100010", 3866 => "10000001", 3868 => "00011000", 3869 => "10110011", 3870 => "00111111", 3871 => "01100011", 3874 => "11000101", 3875 => "00110101", 3877 => "01110001", 3878 => "01101010", 3879 => "10010010", 3880 => "10101000", 3881 => "01100101", 3882 => "10101011", 3883 => "11001110", 3885 => "11001000", 3886 => "01100100", 3889 => "10001000", 3890 => "11100000", 3892 => "11100100", 3893 => "01001111", 3894 => "00101110", 3895 => "11000101", 3896 => "10001001", 3899 => "00101100", 3900 => "00110101", 3903 => "10101000", 3904 => "01000010", 3905 => "10010000", 3906 => "00001000", 3907 => "11110011", 3908 => "11111110", 3909 => "10110011", 3911 => "11100010", 3912 => "00011011", 3913 => "10011101", 3914 => "11101011", 3916 => "10110101", 3917 => "00001010", 3918 => "10011001", 3919 => "01011100", 3920 => "10010010", 3921 => "01010001", 3922 => "10001001", 3923 => "11001011", 3924 => "10111111", 3925 => "11101110", 3927 => "11000101", 3928 => "11111010", 3929 => "11110001", 3930 => "10100000", 3931 => "10001010", 3932 => "00010100", 3933 => "11010011", 3934 => "11100101", 3935 => "01000000", 3937 => "11001011", 3938 => "10011100", 3939 => "10110000", 3941 => "00110100", 3944 => "11011100", 3946 => "11100101", 3947 => "10111100", 3949 => "01101010", 3950 => "01111001", 3951 => "11110011", 3952 => "01000001", 3954 => "01111101", 3956 => "11011101", 3958 => "11001110", 3959 => "00010110", 3961 => "00110001", 3962 => "00100001", 3963 => "10001011", 3964 => "00001000", 3965 => "00000011", 3966 => "11001001", 3967 => "01010010", 3968 => "11011000", 3969 => "01010110", 3970 => "11110000", 3972 => "11100001", 3973 => "11100110", 3975 => "10100101", 3977 => "10110001", 3978 => "10110110", 3979 => "10011100", 3981 => "10000001", 3982 => "01111011", 3983 => "11000110", 3984 => "11000100", 3985 => "11100101", 3986 => "10010000", 3988 => "10110000", 3989 => "10111111", 3990 => "01001010", 3991 => "10111010", 3992 => "10111000", 3993 => "00000110", 3995 => "10010001", 3997 => "11000001", 3998 => "10010000", 3999 => "01100011", 4000 => "01101010", 4001 => "11100111", 4002 => "10001111", 4003 => "10000110", 4004 => "10110110", 4005 => "11010011", 4007 => "01101011", 4008 => "10100000", 4010 => "10101000", 4011 => "11010111", 4012 => "11000011", 4013 => "01101011", 4014 => "11001000", 4015 => "10100001", 4017 => "11011010", 4019 => "11011100", 4020 => "00111011", 4024 => "11011000", 4025 => "10110000", 4026 => "11110001", 4027 => "11010011", 4028 => "01111000", 4029 => "00110101", 4030 => "00110110", 4032 => "00101110", 4033 => "11001010", 4034 => "00100110", 4037 => "10001110", 4038 => "10100001", 4039 => "00110011", 4040 => "10000000", 4044 => "01111101", 4045 => "11010101", 4047 => "00111100", 4048 => "11101001", 4049 => "10001100", 4050 => "00111000", 4052 => "00100100", 4053 => "11110100", 4054 => "10010111", 4055 => "00001110", 4057 => "01010011", 4058 => "01000100", 4059 => "10111001", 4060 => "00011010", 4061 => "01111011", 4062 => "10001010", 4063 => "10100100", 4065 => "01100111", 4067 => "00010001", 4069 => "11101100", 4071 => "00000111", 4074 => "10011111", 4076 => "10100011", 4077 => "01010101", 4080 => "11110000", 4082 => "10111011", 4083 => "11011111", 4087 => "01011010", 4088 => "01011100", 4089 => "00001111", 4090 => "01111010", 4091 => "10111000", 4092 => "01111100", 4094 => "01001011", 4095 => "00010110", 4096 => "10001100", 4097 => "11001011", 4098 => "10111110", 4099 => "10111001", 4100 => "00110100", 4101 => "00001000", 4102 => "01010111", 4106 => "11110111", 4108 => "01001111", 4110 => "10111010", 4111 => "10111011", 4113 => "11101101", 4114 => "01010101", 4115 => "01100110", 4116 => "01010001", 4117 => "01101101", 4118 => "11111011", 4119 => "10111110", 4120 => "01000010", 4121 => "11110000", 4122 => "01010000", 4123 => "01000101", 4124 => "00101100", 4126 => "00100011", 4127 => "11101011", 4128 => "01110001", 4129 => "00011010", 4131 => "11011011", 4132 => "11111000", 4133 => "01011000", 4134 => "11110010", 4135 => "11000010", 4136 => "10000000", 4137 => "10101001", 4139 => "11011000", 4143 => "10110101", 4144 => "00011001", 4145 => "10110000", 4146 => "11100101", 4148 => "11010000", 4149 => "11100011", 4150 => "00101010", 4152 => "01010000", 4154 => "00110100", 4155 => "10110010", 4157 => "01111011", 4158 => "10011000", 4159 => "11011010", 4161 => "11001000", 4162 => "10111111", 4163 => "11000001", 4164 => "11001000", 4165 => "10010011", 4166 => "00110000", 4168 => "10000110", 4169 => "10111101", 4170 => "01011000", 4171 => "00011010", 4173 => "00001011", 4175 => "10111011", 4177 => "10010111", 4178 => "11001101", 4179 => "10110110", 4180 => "01011111", 4181 => "10011011", 4182 => "10110001", 4183 => "10100001", 4184 => "01110001", 4186 => "01011000", 4187 => "01010100", 4188 => "10100101", 4189 => "10100011", 4191 => "10000111", 4192 => "01100110", 4194 => "10100101", 4195 => "10011100", 4196 => "11001111", 4197 => "10101010", 4198 => "00010011", 4199 => "11101110", 4200 => "01000010", 4201 => "10111001", 4202 => "10101100", 4203 => "01100000", 4205 => "10001101", 4207 => "01011011", 4208 => "00110011", 4209 => "01000000", 4211 => "10111111", 4212 => "00001110", 4213 => "00100100", 4214 => "10110000", 4216 => "11111110", 4217 => "11000101", 4218 => "10111110", 4220 => "00001110", 4221 => "11111011", 4222 => "00001011", 4223 => "10011001", 4224 => "10101010", 4225 => "11010011", 4226 => "11100011", 4227 => "11111100", 4228 => "00101001", 4229 => "00101011", 4230 => "01001100", 4232 => "01101101", 4234 => "01000000", 4235 => "01001111", 4236 => "00010111", 4237 => "01101111", 4238 => "11101100", 4239 => "11101010", 4240 => "00110001", 4241 => "11001101", 4242 => "11101010", 4244 => "01000001", 4245 => "11000111", 4246 => "01011100", 4247 => "10100011", 4248 => "01010101", 4250 => "11101111", 4251 => "00010001", 4253 => "00011110", 4254 => "01111011", 4256 => "00111011", 4257 => "00010010", 4258 => "00001000", 4260 => "01110010", 4261 => "00011010", 4263 => "01101111", 4269 => "01100011", 4271 => "11010110", 4272 => "10110001", 4274 => "11111111", 4276 => "01010101", 4280 => "10101100", 4281 => "01011001", 4282 => "10101011", 4283 => "11111101", 4284 => "11110100", 4286 => "01100110", 4288 => "01000000", 4289 => "00101000", 4290 => "00101101", 4291 => "10101101", 4292 => "00010110", 4293 => "01101101", 4294 => "11001001", 4295 => "11001101", 4296 => "00010111", 4301 => "01100001", 4302 => "01000010", 4303 => "10100101", 4305 => "10001000", 4306 => "01000010", 4307 => "10010001", 4309 => "11011000", 4310 => "11010010", 4311 => "00010001", 4312 => "10010100", 4313 => "01000001", 4314 => "11110110", 4315 => "01100011", 4316 => "00001111", 4318 => "01100111", 4319 => "00111011", 4320 => "11010000", 4321 => "00010001", 4323 => "10011100", 4324 => "01000011", 4325 => "11110011", 4326 => "00100111", 4327 => "01001011", 4328 => "10111101", 4330 => "00010111", 4333 => "11010011", 4336 => "01011000", 4337 => "01000110", 4338 => "11001000", 4340 => "10010111", 4341 => "00000110", 4343 => "10000110", 4344 => "00110001", 4345 => "01110011", 4346 => "00010110", 4347 => "11110011", 4348 => "11101011", 4349 => "11000101", 4350 => "11011110", 4351 => "00001010", 4352 => "00110110", 4353 => "10100111", 4354 => "11101100", 4355 => "10011101", 4356 => "01001111", 4357 => "10001001", 4358 => "01001111", 4359 => "01011100", 4360 => "01010001", 4361 => "01100100", 4362 => "10011100", 4363 => "01011010", 4365 => "10000000", 4366 => "10100111", 4367 => "11101000", 4368 => "01110110", 4369 => "10001010", 4370 => "01110010", 4371 => "11110010", 4372 => "11000100", 4373 => "11110100", 4374 => "01011000", 4375 => "00110000", 4377 => "00100001", 4378 => "10110000", 4379 => "11111110", 4380 => "01100000", 4381 => "00001000", 4384 => "01100000", 4387 => "11001110", 4388 => "01001101", 4389 => "11111001", 4390 => "11111101", 4391 => "10110101", 4392 => "00111111", 4393 => "00000110", 4394 => "00010010", 4395 => "11000110", 4397 => "11100100", 4398 => "11000010", 4399 => "01000101", 4402 => "10101010", 4404 => "01101111", 4405 => "00001010", 4406 => "00001010", 4408 => "01101010", 4410 => "11100110", 4411 => "11111101", 4413 => "10101100", 4414 => "00111101", 4415 => "11001101", 4416 => "10010110", 4417 => "01101110", 4418 => "10101100", 4419 => "11011111", 4420 => "00110101", 4424 => "10111110", 4425 => "01011110", 4426 => "11000111", 4429 => "00001000", 4430 => "11110111", 4432 => "01100101", 4433 => "01110001", 4434 => "01001110", 4436 => "00110001", 4437 => "10010011", 4438 => "11001100", 4439 => "10001100", 4440 => "10110010", 4441 => "01000101", 4442 => "11101111", 4444 => "00001001", 4447 => "11101110", 4448 => "01010011", 4449 => "11110001", 4450 => "00001000", 4451 => "00110000", 4452 => "01111100", 4453 => "00111011", 4454 => "00111110", 4456 => "01010101", 4457 => "00111011", 4458 => "10011111", 4459 => "00101010", 4461 => "10000010", 4462 => "01011111", 4463 => "00011010", 4464 => "10011000", 4465 => "01101001", 4467 => "00000101", 4469 => "01111001", 4471 => "00110100", 4472 => "11011100", 4473 => "01100101", 4476 => "00011001", 4477 => "01110100", 4478 => "00111001", 4479 => "11000111", 4480 => "01000011", 4481 => "10010100", 4482 => "01000111", 4483 => "10001110", 4484 => "01110010", 4485 => "10111110", 4486 => "10000111", 4488 => "01101111", 4489 => "01000000", 4490 => "10000011", 4492 => "00100101", 4493 => "10110101", 4495 => "01010010", 4499 => "10011000", 4500 => "01001010", 4501 => "10110111", 4502 => "00001110", 4504 => "00010000", 4505 => "10110000", 4506 => "10010101", 4508 => "00100010", 4509 => "11010110", 4510 => "11000110", 4511 => "00010001", 4513 => "11001110", 4516 => "10110110", 4518 => "01011110", 4519 => "01000001", 4522 => "10010100", 4523 => "11000111", 4524 => "01111010", 4526 => "01010100", 4527 => "10100000", 4528 => "00101001", 4529 => "00010110", 4532 => "00010110", 4533 => "01001100", 4534 => "10010100", 4535 => "01101011", 4536 => "10000101", 4537 => "00010000", 4538 => "10111001", 4539 => "01110011", 4540 => "01101001", 4541 => "01011001", 4543 => "11011110", 4544 => "00101101", 4545 => "01011000", 4546 => "00101010", 4547 => "11000100", 4548 => "01100001", 4549 => "00011001", 4554 => "10101001", 4557 => "00010000", 4558 => "10101000", 4560 => "10101010", 4562 => "11101000", 4563 => "01010110", 4564 => "11011101", 4565 => "11000011", 4566 => "00011111", 4567 => "01100110", 4568 => "10000011", 4570 => "01101101", 4571 => "01101100", 4572 => "11011110", 4573 => "01101110", 4574 => "00000100", 4575 => "10100110", 4576 => "01101111", 4579 => "10001100", 4580 => "11001100", 4582 => "00110111", 4584 => "00100101", 4586 => "00100010", 4587 => "00100101", 4588 => "00010110", 4590 => "10011110", 4594 => "11100001", 4595 => "01001010", 4596 => "00001100", 4597 => "11111010", 4598 => "10000101", 4599 => "00111111", 4600 => "11110100", 4601 => "11111101", 4602 => "01101111", 4604 => "01110001", 4607 => "00100000", 4608 => "01110001", 4612 => "11001000", 4613 => "10001111", 4614 => "11000011", 4615 => "11110111", 4616 => "01110100", 4618 => "01111000", 4619 => "10101011", 4620 => "11100011", 4623 => "01110110", 4624 => "10001101", 4626 => "00110010", 4628 => "10010011", 4629 => "10001111", 4630 => "10001101", 4631 => "00000011", 4632 => "00000011", 4633 => "10100110", 4634 => "10000100", 4638 => "10010000", 4639 => "01100010", 4641 => "10110110", 4642 => "01000001", 4643 => "01011001", 4644 => "11001110", 4646 => "11011100", 4648 => "10001111", 4650 => "11101001", 4651 => "11110010", 4652 => "00010000", 4653 => "10010100", 4654 => "00111001", 4655 => "00101110", 4657 => "00111001", 4658 => "11111010", 4663 => "01100001", 4666 => "01000011", 4668 => "00111100", 4669 => "01000101", 4670 => "00110010", 4671 => "10011000", 4672 => "01100110", 4673 => "11011100", 4674 => "10100000", 4675 => "01100100", 4676 => "00111011", 4677 => "01100010", 4678 => "01110111", 4680 => "01101011", 4681 => "00101010", 4682 => "01100101", 4683 => "01010000", 4684 => "10010000", 4686 => "11100001", 4687 => "11111001", 4688 => "01011100", 4690 => "01110010", 4692 => "10111100", 4694 => "01101110", 4695 => "00000001", 4697 => "10100110", 4699 => "01011001", 4704 => "10101101", 4705 => "00000100", 4706 => "10110011", 4707 => "10101011", 4708 => "01100001", 4709 => "00111110", 4710 => "00000001", 4711 => "10001110", 4713 => "00011110", 4714 => "10010110", 4715 => "01100000", 4716 => "11001000", 4717 => "01001010", 4720 => "11101101", 4721 => "10100111", 4722 => "01000001", 4723 => "10101010", 4726 => "01111011", 4727 => "01111111", 4728 => "01111111", 4729 => "01010100", 4730 => "11101110", 4731 => "10011110", 4736 => "00111101", 4738 => "11011001", 4739 => "10000000", 4740 => "11000001", 4742 => "10110101", 4743 => "01101111", 4744 => "11111100", 4745 => "00101101", 4746 => "00001001", 4747 => "00111001", 4748 => "01100101", 4749 => "00010100", 4750 => "01110010", 4751 => "10000000", 4752 => "11011110", 4753 => "00101010", 4754 => "10101101", 4755 => "01111001", 4758 => "11000110", 4760 => "11100100", 4763 => "11010001", 4764 => "00101010", 4765 => "00111101", 4767 => "10100101", 4768 => "00100100", 4769 => "10010001", 4771 => "01001000", 4773 => "10001101", 4775 => "01001010", 4776 => "10000100", 4778 => "10111010", 4779 => "10010111", 4780 => "10011001", 4781 => "11111001", 4782 => "01011001", 4785 => "01101001", 4787 => "01110010", 4788 => "01101101", 4789 => "10010011", 4790 => "10110001", 4791 => "10011110", 4792 => "11011100", 4795 => "01111101", 4796 => "11100111", 4798 => "10010101", 4799 => "10001111", 4802 => "00110000", 4804 => "10010110", 4805 => "01000101", 4810 => "01111001", 4812 => "10111110", 4813 => "11110100", 4814 => "11000100", 4816 => "10000111", 4817 => "10000100", 4818 => "10110100", 4819 => "00111001", 4820 => "00001100", 4821 => "10100100", 4822 => "00001001", 4823 => "01111100", 4824 => "00010100", 4825 => "00011011", 4827 => "10011110", 4828 => "10010101", 4829 => "11101110", 4830 => "10101100", 4831 => "00100001", 4832 => "00011101", 4833 => "10101100", 4834 => "00110010", 4836 => "00011110", 4837 => "11100010", 4838 => "11101000", 4839 => "10101111", 4840 => "11111110", 4841 => "10011000", 4842 => "11001101", 4843 => "01010011", 4844 => "00000111", 4847 => "11111010", 4848 => "10010010", 4849 => "01111100", 4850 => "11010111", 4851 => "00011111", 4852 => "00011100", 4853 => "01110001", 4856 => "11011001", 4857 => "11101111", 4858 => "01101000", 4859 => "11011010", 4860 => "00101111", 4861 => "11001000", 4862 => "11011011", 4863 => "11100001", 4864 => "11111010", 4865 => "10101100", 4870 => "00111001", 4871 => "00110110", 4872 => "01001010", 4873 => "00101110", 4874 => "00100011", 4875 => "01000110", 4879 => "10001000", 4880 => "00000100", 4881 => "11111001", 4884 => "01110000", 4885 => "11100110", 4886 => "01011101", 4887 => "01100111", 4888 => "00010011", 4891 => "01000001", 4892 => "01101010", 4893 => "11010010", 4894 => "01011110", 4895 => "11010111", 4896 => "11110000", 4897 => "10000111", 4898 => "11000100", 4899 => "00000100", 4900 => "00100110", 4901 => "10000011", 4902 => "01101001", 4903 => "01000010", 4904 => "11001101", 4905 => "00110100", 4906 => "11011100", 4907 => "10101110", 4908 => "10111110", 4909 => "11000110", 4911 => "01011011", 4912 => "00001001", 4913 => "01100100", 4914 => "10011000", 4915 => "11010000", 4916 => "00000111", 4919 => "01000010", 4920 => "00110011", 4921 => "00100101", 4922 => "01010110", 4923 => "10100000", 4924 => "10000000", 4925 => "10001011", 4926 => "10011110", 4927 => "10000010", 4928 => "01000001", 4929 => "01100101", 4930 => "00101000", 4932 => "10010001", 4933 => "11101101", 4934 => "00001110", 4935 => "01001010", 4936 => "01001101", 4937 => "10001000", 4939 => "01001010", 4940 => "10100010", 4941 => "01010011", 4942 => "10010011", 4943 => "10110100", 4944 => "01010000", 4945 => "10110111", 4946 => "00001101", 4948 => "00100101", 4949 => "11100100", 4951 => "00011110", 4952 => "11011110", 4954 => "10000100", 4955 => "01100011", 4956 => "10100111", 4957 => "11111101", 4960 => "00011111", 4961 => "01000011", 4962 => "10110111", 4963 => "01010010", 4964 => "11101100", 4965 => "00011100", 4966 => "11000110", 4967 => "11100111", 4969 => "00000011", 4970 => "10001111", 4971 => "01100110", 4972 => "10011010", 4973 => "11001110", 4975 => "00000100", 4977 => "00010110", 4979 => "10000001", 4980 => "01000010", 4981 => "00111000", 4983 => "00101001", 4984 => "00011010", 4985 => "10001111", 4986 => "11001101", 4987 => "11010100", 4988 => "00010001", 4990 => "00111110", 4991 => "01110110", 4992 => "00110100", 4993 => "10001101", 4995 => "11011110", 4996 => "11010110", 4997 => "10011110", 4999 => "00011111", 5000 => "00101010", 5001 => "01011001", 5003 => "00000100", 5004 => "10001100", 5005 => "11111001", 5008 => "10001101", 5009 => "10000010", 5012 => "01011101", 5015 => "11111110", 5016 => "10111010", 5017 => "00010100", 5018 => "01111100", 5021 => "01111010", 5022 => "10111110", 5023 => "11011100", 5025 => "00010111", 5027 => "01100101", 5029 => "00101100", 5030 => "01011100", 5031 => "10001101", 5032 => "01110000", 5033 => "01010101", 5034 => "10101000", 5038 => "10100001", 5039 => "00011010", 5040 => "11000111", 5043 => "00001110", 5044 => "00111001", 5045 => "11011011", 5046 => "00101010", 5047 => "11110110", 5048 => "00100111", 5050 => "01000001", 5055 => "10001000", 5056 => "00101011", 5057 => "00010011", 5058 => "01001000", 5059 => "01001110", 5060 => "01001011", 5061 => "01011011", 5062 => "10001101", 5063 => "01111011", 5067 => "11001111", 5068 => "10101001", 5069 => "11100001", 5070 => "00010011", 5071 => "00111100", 5073 => "10101100", 5074 => "00000110", 5075 => "10110110", 5076 => "01100110", 5079 => "00000111", 5080 => "11101100", 5081 => "01011110", 5082 => "01000010", 5084 => "00110110", 5085 => "11111100", 5088 => "00100101", 5089 => "10111101", 5090 => "01000000", 5091 => "11110111", 5092 => "01010011", 5093 => "11011101", 5095 => "10101111", 5096 => "10111100", 5097 => "00100111", 5099 => "00101001", 5101 => "11010010", 5103 => "11101100", 5104 => "11001100", 5105 => "11011101", 5106 => "00111000", 5107 => "00110001", 5108 => "00011010", 5109 => "00010111", 5110 => "01011000", 5112 => "00001100", 5113 => "00111010", 5114 => "01011000", 5115 => "00101110", 5116 => "01011111", 5117 => "10100110", 5118 => "00011110", 5119 => "01100100", 5120 => "00010110", 5121 => "01010110", 5122 => "00100111", 5123 => "00111111", 5124 => "10101011", 5126 => "10001111", 5129 => "01011101", 5130 => "00111101", 5132 => "00111100", 5133 => "11010000", 5134 => "11000110", 5135 => "01010111", 5136 => "10000111", 5137 => "11100011", 5140 => "00010110", 5141 => "10001101", 5142 => "00110111", 5144 => "10011111", 5145 => "00010000", 5146 => "11111110", 5148 => "01101011", 5149 => "00000100", 5150 => "10001010", 5152 => "11010110", 5156 => "11011011", 5158 => "01000101", 5161 => "00111110", 5163 => "00011101", 5166 => "10101100", 5167 => "00111000", 5168 => "10000110", 5169 => "11001101", 5171 => "01111100", 5172 => "01111110", 5173 => "10001000", 5174 => "11001110", 5178 => "11111101", 5180 => "00101010", 5181 => "10010101", 5182 => "11111011", 5183 => "10101010", 5184 => "10010010", 5185 => "10010010", 5186 => "00010100", 5187 => "10111100", 5190 => "01100001", 5191 => "00000100", 5192 => "11100010", 5193 => "01100111", 5194 => "01001100", 5195 => "00111110", 5198 => "00001100", 5199 => "10011011", 5200 => "00010010", 5201 => "11011000", 5202 => "10101100", 5203 => "00000010", 5204 => "01111101", 5205 => "11000100", 5208 => "10100111", 5210 => "10001100", 5211 => "01111010", 5213 => "00001000", 5215 => "01010011", 5216 => "11011010", 5217 => "11011110", 5219 => "10100000", 5220 => "00111100", 5221 => "01010111", 5222 => "01000011", 5223 => "01011000", 5224 => "00010100", 5225 => "01001001", 5226 => "11110011", 5227 => "00011111", 5228 => "01110011", 5229 => "11011011", 5230 => "11010101", 5231 => "00101110", 5232 => "01100101", 5233 => "11001001", 5234 => "11100001", 5235 => "00011111", 5236 => "01001100", 5237 => "11111110", 5238 => "01010111", 5239 => "01010011", 5240 => "11010000", 5242 => "01100001", 5243 => "00011000", 5244 => "01001000", 5246 => "10111101", 5248 => "10010001", 5250 => "01010011", 5251 => "10011001", 5252 => "00111000", 5253 => "10011000", 5254 => "00011110", 5255 => "00111010", 5256 => "00111010", 5257 => "00001010", 5258 => "00010101", 5259 => "11001110", 5260 => "01111110", 5261 => "10010010", 5262 => "11111110", 5263 => "01101000", 5265 => "10001001", 5266 => "01011101", 5267 => "11110000", 5270 => "11110100", 5271 => "11111110", 5272 => "10111000", 5273 => "10101001", 5274 => "11010111", 5276 => "10011100", 5277 => "11000010", 5280 => "10110111", 5282 => "01011100", 5285 => "10110010", 5286 => "10000011", 5287 => "00101110", 5289 => "00111101", 5291 => "00000001", 5293 => "01010010", 5294 => "11010100", 5295 => "11000111", 5296 => "11101010", 5297 => "01011011", 5298 => "11100011", 5299 => "01000110", 5300 => "01010000", 5302 => "11111011", 5303 => "11101001", 5305 => "00001111", 5307 => "11001101", 5308 => "00111100", 5309 => "10011010", 5315 => "10010110", 5316 => "10011110", 5320 => "10100010", 5322 => "00000001", 5323 => "11011000", 5324 => "00100111", 5325 => "10000100", 5326 => "10011001", 5327 => "00010010", 5328 => "11000110", 5329 => "11010101", 5332 => "00110101", 5333 => "00011011", 5335 => "01100011", 5336 => "00101101", 5337 => "11000101", 5338 => "00010011", 5339 => "11010011", 5340 => "00010100", 5341 => "01110111", 5342 => "10000000", 5343 => "01101100", 5345 => "11000110", 5346 => "01000100", 5347 => "11001111", 5349 => "00001000", 5350 => "11001110", 5351 => "01110010", 5352 => "01101100", 5353 => "01001001", 5354 => "11100010", 5355 => "10111001", 5356 => "01110111", 5357 => "11011111", 5358 => "00101010", 5359 => "11001101", 5360 => "00000011", 5361 => "00111110", 5363 => "00011010", 5364 => "11111011", 5365 => "01000000", 5367 => "01100111", 5368 => "11110100", 5370 => "01001011", 5373 => "00100110", 5374 => "10010101", 5377 => "10100000", 5378 => "10010001", 5379 => "11101011", 5380 => "11011110", 5382 => "10010101", 5383 => "01011100", 5385 => "00100111", 5387 => "01001110", 5388 => "10000110", 5389 => "10001110", 5391 => "11011111", 5393 => "01010001", 5394 => "00011011", 5395 => "11011100", 5397 => "00110001", 5398 => "00001111", 5399 => "00101011", 5401 => "01110101", 5403 => "10011101", 5404 => "10010011", 5406 => "11000101", 5407 => "10010111", 5408 => "00100110", 5411 => "10010110", 5412 => "01001111", 5413 => "01100000", 5414 => "11010001", 5415 => "01001110", 5416 => "10010110", 5417 => "11000101", 5419 => "11100011", 5420 => "01100001", 5422 => "11010100", 5424 => "00100000", 5425 => "01111011", 5426 => "10000001", 5427 => "01101111", 5428 => "11110000", 5429 => "11101010", 5430 => "10010100", 5431 => "00001100", 5432 => "10111000", 5433 => "11010001", 5434 => "01000101", 5436 => "01101100", 5437 => "10111100", 5438 => "10101001", 5440 => "00011100", 5442 => "11010001", 5444 => "01001101", 5446 => "11011101", 5448 => "11111010", 5449 => "01011100", 5450 => "11001010", 5451 => "00110111", 5452 => "01100011", 5453 => "00011101", 5455 => "00011000", 5457 => "01111011", 5458 => "11100100", 5459 => "11000010", 5460 => "10010101", 5462 => "10010000", 5463 => "10001100", 5464 => "10101010", 5466 => "11110011", 5468 => "01101001", 5469 => "01101000", 5471 => "10001011", 5472 => "11000010", 5473 => "11011100", 5474 => "00100010", 5475 => "01000101", 5476 => "01010111", 5478 => "11001011", 5479 => "01110001", 5480 => "11100001", 5483 => "10010111", 5486 => "01100110", 5488 => "11001111", 5489 => "00000011", 5490 => "11101000", 5491 => "00001000", 5493 => "11100011", 5494 => "00101100", 5496 => "10111101", 5498 => "01110011", 5499 => "00011010", 5500 => "01101101", 5502 => "11010011", 5503 => "01111100", 5504 => "11001100", 5506 => "01110010", 5507 => "10011100", 5509 => "10101100", 5510 => "01100011", 5511 => "11110001", 5512 => "11010000", 5513 => "10011100", 5514 => "01011110", 5516 => "10111111", 5517 => "00011001", 5518 => "11110110", 5519 => "01100011", 5520 => "10101010", 5521 => "10000101", 5522 => "01111101", 5525 => "01111010", 5526 => "00101110", 5527 => "11011100", 5529 => "00001111", 5530 => "00010101", 5531 => "11000110", 5532 => "10011101", 5533 => "01000010", 5534 => "11000111", 5535 => "11010011", 5536 => "01010001", 5537 => "10001010", 5538 => "10001000", 5540 => "00011011", 5541 => "01011100", 5542 => "10000000", 5543 => "10010111", 5544 => "10111101", 5545 => "11100001", 5546 => "11001011", 5547 => "00100111", 5548 => "10000000", 5550 => "11000111", 5552 => "10011111", 5553 => "11010011", 5554 => "01001010", 5555 => "01000001", 5556 => "11000000", 5557 => "10101111", 5558 => "11111011", 5559 => "11011011", 5560 => "01101100", 5561 => "10010010", 5562 => "10110100", 5563 => "11100110", 5564 => "01100111", 5565 => "11110110", 5566 => "11000010", 5569 => "10010100", 5570 => "01010111", 5571 => "01000011", 5572 => "00100100", 5573 => "00010100", 5574 => "11100000", 5576 => "00101000", 5577 => "10101001", 5578 => "11101100", 5579 => "01110111", 5580 => "01001100", 5585 => "11101111", 5586 => "10010110", 5587 => "10100010", 5588 => "01100111", 5590 => "01010001", 5591 => "01000110", 5592 => "11110100", 5593 => "10001000", 5596 => "11011101", 5598 => "10001000", 5599 => "01100101", 5600 => "00001001", 5601 => "00111011", 5602 => "10111100", 5603 => "01110110", 5604 => "11010100", 5605 => "10110010", 5606 => "00101100", 5607 => "10001001", 5608 => "11100001", 5609 => "01110001", 5610 => "11000010", 5611 => "11000001", 5612 => "01101000", 5613 => "10101001", 5614 => "01001110", 5615 => "00000011", 5616 => "01000100", 5617 => "00101011", 5618 => "01110111", 5619 => "10110011", 5622 => "01111101", 5623 => "01001110", 5625 => "01010010", 5627 => "00010110", 5628 => "10000000", 5630 => "00101010", 5632 => "00010010", 5634 => "11110000", 5635 => "11101011", 5636 => "10101011", 5637 => "11101101", 5639 => "10001010", 5641 => "00001101", 5643 => "00000011", 5644 => "01111100", 5645 => "11000101", 5646 => "01111101", 5648 => "10101010", 5649 => "11110100", 5652 => "00100110", 5653 => "00111010", 5655 => "00011100", 5656 => "11000010", 5657 => "11011000", 5658 => "10001100", 5660 => "11101110", 5661 => "00010010", 5662 => "01001111", 5664 => "11110101", 5665 => "01100100", 5666 => "01111011", 5667 => "00010110", 5668 => "11110001", 5670 => "10011101", 5671 => "10010111", 5672 => "01101011", 5673 => "01111011", 5675 => "10101110", 5677 => "11101100", 5678 => "01001010", 5679 => "01100011", 5680 => "10110001", 5681 => "10011001", 5685 => "11000100", 5686 => "11000010", 5687 => "01100100", 5688 => "11001100", 5693 => "01101000", 5694 => "10101101", 5697 => "10110110", 5698 => "10001111", 5699 => "10110001", 5702 => "11100000", 5703 => "10100011", 5704 => "01001010", 5706 => "01001100", 5707 => "10000101", 5708 => "11101100", 5709 => "00010000", 5710 => "10101000", 5713 => "11110111", 5714 => "10010000", 5715 => "10101101", 5718 => "10001010", 5721 => "10110110", 5722 => "11000011", 5724 => "11101010", 5725 => "10111100", 5727 => "11100101", 5728 => "01011101", 5730 => "00000111", 5731 => "00101001", 5732 => "01001001", 5733 => "00110110", 5734 => "11100111", 5735 => "01001000", 5736 => "01111001", 5737 => "01101110", 5738 => "01110010", 5740 => "11011111", 5741 => "01010000", 5742 => "10000111", 5743 => "00011101", 5744 => "00100111", 5745 => "10110010", 5746 => "01000110", 5747 => "10010001", 5748 => "11001100", 5749 => "00000110", 5751 => "00100111", 5753 => "10110011", 5755 => "11010101", 5756 => "00001010", 5757 => "00111110", 5758 => "00110010", 5759 => "01010010", 5760 => "10010110", 5761 => "11110011", 5762 => "00000010", 5763 => "10101000", 5764 => "10101111", 5765 => "11001101", 5766 => "11111110", 5767 => "11010011", 5768 => "01101111", 5769 => "01000110", 5770 => "10100101", 5771 => "10001111", 5772 => "00111101", 5773 => "01101000", 5774 => "10100010", 5777 => "11110001", 5778 => "11101010", 5779 => "10001010", 5780 => "01111011", 5782 => "10101001", 5783 => "10001010", 5784 => "00010011", 5785 => "10111000", 5786 => "00000111", 5787 => "10110010", 5788 => "10100011", 5790 => "10111100", 5791 => "01000110", 5792 => "01010101", 5793 => "10000000", 5794 => "10010000", 5795 => "11001101", 5797 => "10000000", 5798 => "00110011", 5799 => "01001010", 5801 => "10000110", 5802 => "10011001", 5803 => "00111010", 5804 => "01101100", 5805 => "11001110", 5806 => "00100000", 5807 => "10001000", 5809 => "11001001", 5811 => "01111001", 5812 => "01110001", 5814 => "01111101", 5815 => "00101101", 5816 => "01111010", 5817 => "11001100", 5819 => "00011011", 5821 => "01001000", 5823 => "11110101", 5824 => "00011010", 5825 => "00000110", 5826 => "11011100", 5827 => "10101100", 5829 => "01000011", 5830 => "10100110", 5831 => "11000101", 5832 => "10110110", 5833 => "01010101", 5834 => "00110100", 5835 => "00101000", 5836 => "10011010", 5837 => "11001000", 5838 => "00110100", 5839 => "11111011", 5840 => "10000001", 5841 => "10100101", 5843 => "00010101", 5844 => "00101010", 5845 => "10110011", 5846 => "11101110", 5847 => "10100001", 5848 => "00101111", 5849 => "10001001", 5850 => "10010001", 5851 => "01111011", 5853 => "11101110", 5854 => "01001111", 5855 => "00001000", 5856 => "10111001", 5857 => "11100100", 5858 => "00101010", 5860 => "10011001", 5861 => "10100111", 5871 => "10100110", 5873 => "01001100", 5875 => "11110101", 5877 => "00111000", 5880 => "11010010", 5881 => "01000000", 5882 => "10010100", 5885 => "11001000", 5887 => "10110111", 5888 => "10010110", 5889 => "01111001", 5890 => "11000101", 5891 => "11110110", 5892 => "11000000", 5894 => "10111110", 5895 => "01101011", 5897 => "01100110", 5900 => "01011000", 5901 => "11000001", 5906 => "01110010", 5907 => "10011010", 5909 => "01001110", 5910 => "01111010", 5914 => "00000101", 5915 => "11111111", 5918 => "10001010", 5919 => "11001101", 5921 => "10101111", 5923 => "11100010", 5924 => "00001010", 5925 => "11101111", 5926 => "10110111", 5927 => "00101101", 5928 => "10001110", 5929 => "10000011", 5930 => "11101010", 5931 => "00101001", 5933 => "10010101", 5935 => "00110100", 5936 => "11011010", 5938 => "10110101", 5940 => "00001001", 5941 => "10111110", 5945 => "01001010", 5952 => "11101011", 5955 => "10110100", 5956 => "11111000", 5958 => "00111111", 5959 => "11100011", 5960 => "01010010", 5961 => "10010010", 5963 => "11011111", 5966 => "10101111", 5969 => "10110111", 5970 => "11001000", 5972 => "11000001", 5974 => "11110001", 5976 => "00100110", 5977 => "11011011", 5979 => "11010100", 5980 => "11100110", 5981 => "01101000", 5982 => "00000101", 5983 => "00010111", 5984 => "11110000", 5987 => "00001101", 5988 => "01001000", 5989 => "11110100", 5990 => "00001101", 5991 => "10101001", 5992 => "00010110", 5998 => "10111111", 6000 => "00101110", 6003 => "01100101", 6004 => "01110010", 6005 => "11111111", 6007 => "11101011", 6008 => "11100101", 6010 => "00111001", 6011 => "11111110", 6012 => "10010111", 6014 => "11001100", 6016 => "10000011", 6017 => "11010010", 6018 => "10011101", 6019 => "11001111", 6020 => "01011101", 6023 => "00000110", 6024 => "01111101", 6027 => "11101001", 6029 => "10100011", 6030 => "00110110", 6035 => "11001010", 6036 => "01011101", 6041 => "01110100", 6043 => "11110010", 6045 => "11000001", 6047 => "10101001", 6049 => "10010111", 6050 => "00010000", 6053 => "01100111", 6054 => "10011011", 6056 => "10111100", 6057 => "11010011", 6060 => "00100101", 6066 => "10001110", 6067 => "10011110", 6068 => "11111111", 6069 => "10111111", 6071 => "10010001", 6072 => "00011000", 6074 => "00000100", 6075 => "00100010", 6076 => "00100110", 6078 => "11111110", 6080 => "01000111", 6082 => "01010011", 6083 => "00011010", 6084 => "01000011", 6088 => "01001001", 6089 => "01111111", 6091 => "11100001", 6093 => "00000011", 6096 => "11011100", 6103 => "01001110", 6104 => "10110011", 6105 => "01011000", 6107 => "11001000", 6108 => "01101010", 6110 => "00011000", 6111 => "00101000", 6113 => "00111111", 6114 => "10111011", 6119 => "10110101", 6120 => "01000010", 6123 => "00001101", 6124 => "10010101", 6125 => "10001011", 6127 => "01000100", 6136 => "10001101", 6137 => "11011010", 6138 => "00011000", 6139 => "00010111", 6142 => "11010010", 6143 => "11010011", 6145 => "00010110", 6147 => "10111110", 6149 => "11110001", 6150 => "11000010", 6151 => "10110110", 6152 => "00110001", 6154 => "10010011", 6155 => "10110111", 6157 => "01101100", 6159 => "01110100", 6160 => "11110010", 6162 => "01001101", 6163 => "11000010", 6164 => "10001010", 6165 => "11101110", 6166 => "10100011", 6168 => "00101011", 6169 => "01100110", 6170 => "01011101", 6172 => "01111001", 6173 => "10101100", 6175 => "10111000", 6177 => "10101011", 6185 => "00101110", 6188 => "00110001", 6189 => "11011110", 6191 => "11010000", 6194 => "01010101", 6195 => "01011000", 6196 => "00100010", 6197 => "11010000", 6200 => "00101101", 6202 => "11101001", 6203 => "00100000", 6205 => "11011011", 6207 => "00111101", 6208 => "10011011", 6210 => "11100001", 6213 => "01011001", 6216 => "11010110", 6218 => "01001011", 6220 => "11101010", 6223 => "11100101", 6225 => "01011001", 6228 => "11101000", 6230 => "11100001", 6233 => "11101000", 6234 => "10111100", 6238 => "10101001", 6241 => "00011001", 6247 => "00010011", 6248 => "00100111", 6251 => "10010111", 6253 => "10011101", 6254 => "10010011", 6255 => "01001100", 6256 => "11100100", 6257 => "00010010", 6258 => "11100110", 6260 => "10011110", 6262 => "00100000", 6265 => "10010000", 6266 => "11110001", 6271 => "00010100", 6274 => "01100000", 6275 => "11010000", 6278 => "01000010", 6280 => "00000100", 6282 => "00101101", 6284 => "11011111", 6287 => "11000111", 6288 => "00110111", 6290 => "11111011", 6292 => "00111001", 6294 => "11001000", 6297 => "01101011", 6298 => "10000010", 6302 => "00101111", 6303 => "11001110", 6304 => "11100001", 6305 => "11110100", 6307 => "10000100", 6310 => "10110101", 6312 => "10000110", 6314 => "11111100", 6317 => "11111000", 6319 => "10101100", 6321 => "00101001", 6323 => "11011101", 6326 => "10100101", 6336 => "01111001", 6341 => "10011000", 6344 => "10100000", 6345 => "11101101", 6346 => "01011110", 6347 => "11111111", 6351 => "10100110", 6352 => "11001011", 6356 => "10100110", 6358 => "11011100", 6359 => "00001110", 6360 => "01010110", 6366 => "00110110", 6367 => "11111110", 6369 => "01011101", 6370 => "00001110", 6372 => "10100111", 6373 => "01100111", 6374 => "00001010", 6376 => "00110111", 6377 => "00010100", 6378 => "10101000", 6379 => "00100011", 6380 => "00010100", 6381 => "11001001", 6383 => "00111111", 6387 => "10010011", 6388 => "11010110", 6389 => "00011111", 6392 => "00110011", 6395 => "11001111", 6398 => "01011100", 6400 => "11100000", 6403 => "00100111", 6405 => "11011010", 6411 => "11010100", 6412 => "11111000", 6417 => "00001001", 6419 => "01110101", 6421 => "11011011", 6424 => "11011011", 6425 => "10110100", 6426 => "00000010", 6427 => "00011111", 6428 => "11001100", 6430 => "10100001", 6431 => "11111010", 6436 => "01001011", 6437 => "00011010", 6438 => "00111100", 6441 => "00101011", 6444 => "11010000", 6447 => "11001111", 6448 => "00111111", 6449 => "01000100", 6452 => "00110011", 6456 => "00000100", 6458 => "11001011", 6460 => "01011100", 6462 => "01011101", 6463 => "00010000", 6464 => "01010111", 6465 => "00010011", 6467 => "00110101", 6468 => "01101010", 6469 => "11110110", 6470 => "10111111", 6472 => "10111001", 6475 => "01111010", 6476 => "00100001", 6477 => "01001011", 6479 => "00010010", 6482 => "01010001", 6484 => "10001110", 6486 => "00111111", 6488 => "10100111", 6491 => "01110011", 6493 => "01011101", 6499 => "11100000", 6504 => "00111000", 6505 => "01111110", 6507 => "01000001", 6509 => "10010100", 6511 => "10000110", 6514 => "00101110", 6515 => "00010100", 6522 => "11010111", 6524 => "10000001", 6526 => "11111100", 6527 => "11000000", 6528 => "10110110", 6530 => "11101110", 6533 => "00111100", 6534 => "00010011", 6535 => "10011011", 6537 => "01011101", 6539 => "00100111", 6542 => "10111011", 6545 => "10110110", 6546 => "11001111", 6547 => "01001101", 6548 => "11011100", 6550 => "01010111", 6554 => "00110110", 6555 => "11011101", 6557 => "10001000", 6558 => "10110110", 6561 => "00001001", 6564 => "10001000", 6568 => "00100001", 6570 => "01011000", 6571 => "01001010", 6573 => "01000011", 6575 => "11001001", 6577 => "11001011", 6579 => "10000100", 6580 => "00011101", 6581 => "10001110", 6582 => "00001100", 6583 => "01000010", 6584 => "10001111", 6587 => "10110000", 6588 => "00011111", 6590 => "01000100", 6591 => "00111000", 6593 => "01100100", 6598 => "10101001", 6599 => "11011010", 6601 => "01001110", 6602 => "11010101", 6603 => "00100001", 6605 => "01000010", 6608 => "00000110", 6613 => "00110101", 6614 => "01111101", 6615 => "01101010", 6616 => "01001011", 6617 => "11000011", 6618 => "10101110", 6624 => "10001001", 6626 => "01010010", 6628 => "10011111", 6631 => "10110110", 6633 => "10100111", 6634 => "00011101", 6635 => "00110011", 6637 => "11100001", 6641 => "00000111", 6644 => "01111111", 6645 => "00100111", 6647 => "00101000", 6648 => "11100101", 6649 => "10011111", 6650 => "11000111", 6652 => "10101110", 6656 => "10010001", 6657 => "01000100", 6659 => "00011010", 6660 => "11010111", 6661 => "00000101", 6662 => "00110111", 6663 => "00001110", 6665 => "01100010", 6669 => "10110110", 6670 => "00001111", 6671 => "01100000", 6673 => "01100100", 6675 => "00011110", 6685 => "11011101", 6686 => "10111100", 6688 => "11000110", 6690 => "01101101", 6691 => "01011000", 6694 => "01101001", 6695 => "11010110", 6698 => "01110100", 6699 => "00101010", 6701 => "10101001", 6703 => "00101011", 6704 => "10101101", 6705 => "01010011", 6706 => "11111110", 6707 => "00011001", 6710 => "00001100", 6711 => "00100010", 6712 => "11000010", 6713 => "10001110", 6715 => "10101111", 6718 => "01011110", 6720 => "10110101", 6726 => "00100101", 6727 => "00001100", 6731 => "11000011", 6733 => "00110000", 6736 => "00011011", 6738 => "01110101", 6744 => "01001100", 6746 => "11000010", 6747 => "01111000", 6757 => "00010011", 6761 => "10001110", 6762 => "01011011", 6763 => "01110001", 6765 => "10011000", 6767 => "00001001", 6771 => "10111110", 6772 => "10011110", 6773 => "01001011", 6775 => "10111011", 6776 => "00000111", 6779 => "11100001", 6781 => "00101010", 6783 => "11011010", 6784 => "01001111", 6788 => "10101100", 6792 => "01111010", 6793 => "10011010", 6797 => "01011001", 6799 => "00100001", 6800 => "10001001", 6803 => "10100010", 6806 => "00111101", 6810 => "01101000", 6811 => "10101001", 6815 => "10001011", 6817 => "10001001", 6818 => "10011111", 6820 => "01110010", 6821 => "00101000", 6823 => "01000000", 6824 => "11101000", 6831 => "11000011", 6832 => "01001000", 6834 => "10110100", 6835 => "11000010", 6839 => "11000000", 6840 => "00000001", 6842 => "11101100", 6844 => "11001011", 6845 => "00111111", 6850 => "10101011", 6851 => "11111100", 6855 => "01001010", 6856 => "11111010", 6859 => "11010110", 6860 => "01000010", 6861 => "01111010", 6863 => "01000110", 6864 => "01011001", 6865 => "10011100", 6873 => "00001111", 6874 => "10110001", 6875 => "10001101", 6877 => "10110101", 6879 => "10110100", 6880 => "11111010", 6883 => "00001011", 6884 => "11010111", 6885 => "01111000", 6889 => "01001100", 6898 => "10000010", 6900 => "11101101", 6902 => "00111011", 6903 => "10010000", 6905 => "10110111", 6906 => "01110010", 6908 => "00100101", 6910 => "01100011", 6911 => "01101111", 6914 => "00111100", 6917 => "00100100", 6922 => "00111010", 6923 => "00010011", 6924 => "11000000", 6926 => "10011000", 6928 => "11101010", 6929 => "10101100", 6930 => "11010011", 6933 => "00111101", 6936 => "10110110", 6940 => "11001101", 6941 => "11001010", 6949 => "01010001", 6950 => "10001100", 6952 => "11101010", 6954 => "11111100", 6956 => "10101001", 6957 => "11000000", 6958 => "10110111", 6961 => "01001000", 6962 => "00000101", 6968 => "00010111", 6974 => "00100110", 6978 => "10111100", 6980 => "10001111", 6981 => "00000111", 6983 => "10001100", 6984 => "10111100", 6985 => "10111001", 6988 => "00011011", 6989 => "10001100", 6991 => "10001000", 6993 => "10010010", 6995 => "11101001", 6996 => "11000001", 6998 => "00101001", 7004 => "00101110", 7007 => "11111000", 7008 => "01111110", 7009 => "00100000", 7010 => "11100100", 7015 => "00001110", 7018 => "01011011", 7019 => "11100000", 7020 => "10001010", 7021 => "01100000", 7024 => "01000000", 7025 => "11001100", 7026 => "01010011", 7027 => "01101111", 7028 => "01011111", 7032 => "10010101", 7034 => "11101000", 7035 => "10011001", 7036 => "00011000", 7040 => "00100100", 7045 => "00100110", 7046 => "01100000", 7047 => "10110111", 7048 => "10101111", 7050 => "01010000", 7055 => "10011110", 7058 => "00101011", 7061 => "10011101", 7062 => "01000011", 7063 => "00100101", 7064 => "10110001", 7066 => "00011111", 7067 => "01110010", 7075 => "11110100", 7076 => "00101011", 7077 => "01000011", 7080 => "01000011", 7081 => "10000100", 7086 => "10001001", 7088 => "00100001", 7089 => "01000100", 7090 => "01111111", 7091 => "11001011", 7099 => "10111000", 7100 => "00000100", 7102 => "00010101", 7104 => "00010011", 7106 => "00111101", 7108 => "10101100", 7109 => "00100100", 7110 => "10100010", 7114 => "10000001", 7115 => "10010000", 7116 => "01000111", 7117 => "01111110", 7118 => "10100011", 7122 => "10110110", 7126 => "01100001", 7128 => "11001111", 7129 => "01011011", 7130 => "10011101", 7133 => "00100101", 7134 => "00111101", 7136 => "00101010", 7137 => "10001110", 7138 => "01010101", 7139 => "01011000", 7141 => "01101110", 7142 => "01110001", 7143 => "10101010", 7145 => "01100110", 7148 => "11000111", 7151 => "00100100", 7153 => "10010010", 7154 => "00110110", 7156 => "10101011", 7159 => "01010010", 7163 => "10011111", 7164 => "11111100", 7171 => "10010010", 7173 => "11101011", 7174 => "01100110", 7175 => "10011110", 7177 => "01110111", 7181 => "00111000", 7182 => "10101001", 7187 => "01000011", 7188 => "10110000", 7190 => "00111100", 7193 => "11100000", 7194 => "00000101", 7196 => "00101001", 7200 => "10010001", 7201 => "10101100", 7202 => "01111111", 7203 => "11111011", 7204 => "11001010", 7206 => "10100100", 7208 => "11001110", 7209 => "11000110", 7210 => "10101101", 7212 => "10111100", 7214 => "01011011", 7217 => "01110111", 7219 => "10001101", 7221 => "01100101", 7223 => "11111100", 7227 => "11000010", 7228 => "00110100", 7230 => "01001010", 7232 => "11110111", 7234 => "10010001", 7236 => "11101101", 7237 => "10011000", 7238 => "01100011", 7239 => "01101110", 7242 => "11010000", 7245 => "10000110", 7246 => "11001010", 7250 => "10010010", 7252 => "01100100", 7253 => "10010100", 7254 => "10111101", 7255 => "00101100", 7256 => "00001101", 7260 => "00010101", 7262 => "10010110", 7267 => "10111000", 7268 => "11110010", 7269 => "10010000", 7270 => "01000011", 7272 => "11000010", 7273 => "01110011", 7274 => "01001100", 7279 => "01111111", 7280 => "10110110", 7282 => "10111111", 7286 => "01100111", 7287 => "11101111", 7291 => "10000010", 7295 => "11011111", 7297 => "10011011", 7300 => "00000101", 7302 => "00010001", 7303 => "10100011", 7304 => "00110011", 7308 => "01110011", 7309 => "10111010", 7310 => "00011011", 7313 => "10101001", 7321 => "10010000", 7322 => "00101000", 7326 => "00110010", 7328 => "10010110", 7329 => "01001011", 7331 => "10111101", 7337 => "10011101", 7338 => "00000011", 7339 => "01000011", 7340 => "01001110", 7342 => "00010111", 7345 => "10011110", 7346 => "00011100", 7347 => "11100011", 7351 => "10010100", 7353 => "00011100", 7357 => "01001101", 7361 => "00110011", 7362 => "01101001", 7363 => "00110011", 7364 => "10010001", 7365 => "11000001", 7367 => "00010001", 7368 => "01000011", 7373 => "11000100", 7374 => "00000010", 7375 => "11001000", 7378 => "11100001", 7385 => "11011011", 7388 => "00111100", 7390 => "01101000", 7392 => "01011010", 7393 => "11101101", 7395 => "10110000", 7396 => "01010100", 7400 => "11001101", 7401 => "10100110", 7402 => "00101111", 7403 => "10100000", 7404 => "10010001", 7406 => "10100101", 7409 => "01010011", 7414 => "00100001", 7415 => "01010001", 7422 => "01110011", 7423 => "11011110", 7424 => "01100100", 7426 => "01010111", 7427 => "00011000", 7428 => "01100001", 7430 => "01111010", 7433 => "11101000", 7434 => "11001100", 7436 => "01001010", 7448 => "10000011", 7450 => "11010110", 7453 => "10000010", 7457 => "00011000", 7460 => "11111111", 7461 => "01110101", 7462 => "01011100", 7464 => "11100110", 7465 => "11100100", 7466 => "01101100", 7467 => "01101100", 7469 => "00101100", 7470 => "10100011", 7474 => "10111111", 7475 => "00000110", 7476 => "10001011", 7478 => "10111010", 7480 => "00011001", 7481 => "01110011", 7482 => "11111010", 7483 => "00110011", 7486 => "10101010", 7487 => "10100000", 7488 => "01000101", 7489 => "10111101", 7490 => "01110011", 7497 => "11000111", 7498 => "00010100", 7499 => "10111111", 7500 => "00001010", 7502 => "00000001", 7504 => "00100011", 7505 => "10100111", 7507 => "00100101", 7509 => "10010011", 7510 => "10011111", 7511 => "01111010", 7513 => "00110100", 7514 => "00010000", 7515 => "00101001", 7518 => "11100000", 7519 => "10111001", 7521 => "10000101", 7523 => "01011101", 7524 => "00000101", 7525 => "00110100", 7526 => "00111011", 7527 => "00000001", 7529 => "11111010", 7532 => "00111010", 7534 => "11011111", 7535 => "00111000", 7537 => "11000011", 7538 => "10101101", 7544 => "00000001", 7545 => "10100100", 7547 => "00001111", 7550 => "01110011", 7551 => "01011111", 7552 => "00010110", 7553 => "10010100", 7554 => "01110001", 7557 => "10000110", 7562 => "01111110", 7563 => "11101001", 7567 => "00010100", 7568 => "11001110", 7573 => "10001001", 7576 => "10111000", 7578 => "11011111", 7579 => "11111011", 7580 => "00010000", 7582 => "00100001", 7587 => "11010100", 7589 => "10001011", 7590 => "11111010", 7591 => "11101110", 7596 => "11110001", 7597 => "11110001", 7599 => "00000101", 7601 => "11100110", 7602 => "00101000", 7603 => "00100010", 7604 => "00100000", 7605 => "01010100", 7606 => "00001100", 7608 => "10101101", 7611 => "11010100", 7612 => "10000011", 7619 => "10111110", 7621 => "00011100", 7630 => "10011101", 7634 => "01101010", 7638 => "10011000", 7640 => "01111011", 7644 => "01011101", 7646 => "00001101", 7647 => "00110110", 7654 => "11101000", 7659 => "00011100", 7660 => "11111101", 7661 => "11110011", 7665 => "00010110", 7669 => "10101101", 7670 => "01000000", 7673 => "10001011", 7674 => "10101110", 7676 => "10111011", 7678 => "00001000", 7679 => "10000001", 7681 => "00101111", 7682 => "00000101", 7684 => "11011100", 7685 => "11011110", 7686 => "00110001", 7691 => "11011010", 7694 => "10100110", 7696 => "10010100", 7699 => "00010111", 7700 => "11111010", 7702 => "00011100", 7706 => "10100011", 7707 => "01100000", 7710 => "10001110", 7711 => "10001001", 7717 => "10110101", 7720 => "10011111", 7721 => "00011111", 7723 => "10001110", 7725 => "11110010", 7727 => "01101100", 7728 => "11100000", 7730 => "01001100", 7731 => "01101000", 7733 => "11000100", 7739 => "11110100", 7741 => "11011110", 7744 => "00000011", 7747 => "10010010", 7749 => "00101001", 7754 => "11101001", 7755 => "00100111", 7756 => "01011100", 7757 => "00111000", 7758 => "01100000", 7759 => "00101001", 7760 => "11011111", 7762 => "11100101", 7763 => "11011000", 7764 => "00001010", 7765 => "01010001", 7766 => "10010001", 7767 => "01101100", 7768 => "00111101", 7771 => "01111001", 7774 => "10101000", 7779 => "11100011", 7780 => "11001010", 7783 => "10001101", 7784 => "01100001", 7787 => "10010101", 7790 => "10010110", 7792 => "10000001", 7796 => "11010111", 7798 => "11111001", 7802 => "11001000", 7804 => "11011001", 7805 => "00001100", 7806 => "11010110", 7807 => "11101000", 7811 => "01100111", 7812 => "11011111", 7814 => "01100011", 7818 => "01100100", 7825 => "00100010", 7826 => "10010000", 7827 => "10101010", 7832 => "01110110", 7835 => "10001000", 7836 => "01001111", 7839 => "10101011", 7840 => "11100000", 7843 => "01011110", 7846 => "10101001", 7847 => "01110111", 7848 => "11101001", 7850 => "00100111", 7853 => "00100101", 7854 => "01010010", 7855 => "10010101", 7856 => "11100110", 7857 => "00001110", 7859 => "00100111", 7860 => "10011110", 7862 => "00101010", 7864 => "00000001", 7866 => "11101111", 7869 => "00100101", 7870 => "10010101", 7871 => "11100100", 7873 => "11111110", 7877 => "11011111", 7879 => "10011100", 7885 => "01111110", 7886 => "00001110", 7887 => "01100000", 7888 => "01100010", 7889 => "11001011", 7891 => "11111010", 7895 => "00111110", 7897 => "01001010", 7899 => "01010100", 7900 => "10011100", 7904 => "11110111", 7907 => "01111100", 7910 => "10101101", 7915 => "10001001", 7916 => "00001000", 7918 => "00010110", 7919 => "01010101", 7920 => "01100101", 7921 => "11010011", 7923 => "10000010", 7924 => "01100010", 7926 => "00100111", 7927 => "01111001", 7930 => "00010100", 7932 => "11011101", 7933 => "01011110", 7935 => "10111101", 7936 => "11001110", 7940 => "10110000", 7941 => "10000100", 7945 => "01100110", 7946 => "00000010", 7947 => "10001011", 7950 => "11000001", 7951 => "01010001", 7953 => "01101000", 7954 => "10110100", 7955 => "10011101", 7956 => "11010000", 7957 => "10011011", 7959 => "11110100", 7966 => "00100101", 7967 => "00110000", 7970 => "01110110", 7971 => "00110010", 7972 => "10111100", 7973 => "00011001", 7976 => "01011000", 7979 => "01101100", 7980 => "11100010", 7982 => "00011100", 7983 => "11010010", 7984 => "00001100", 7986 => "10101101", 7988 => "11000011", 7990 => "01110100", 7991 => "10100010", 7992 => "10000100", 7994 => "01100000", 7997 => "01001101", 7998 => "00100101", 8003 => "00100100", 8004 => "11001011", 8005 => "00010110", 8006 => "01000110", 8008 => "01010001", 8009 => "10111110", 8010 => "00100001", 8011 => "01000111", 8013 => "11111110", 8015 => "11101011", 8017 => "00100111", 8018 => "11110011", 8019 => "00011010", 8025 => "00101110", 8030 => "00011010", 8033 => "11001010", 8034 => "11000011", 8036 => "01110110", 8037 => "11001110", 8038 => "11010010", 8041 => "01010011", 8042 => "11100001", 8044 => "01110110", 8045 => "11000010", 8048 => "10110000", 8052 => "11111110", 8053 => "11000001", 8054 => "00100100", 8055 => "10110101", 8057 => "10111110", 8059 => "11100101", 8062 => "11010010", 8066 => "01011100", 8067 => "11110000", 8068 => "10001000", 8069 => "00111110", 8073 => "11110110", 8074 => "11000101", 8075 => "01010110", 8079 => "01001010", 8087 => "10110101", 8090 => "00101110", 8091 => "10110100", 8092 => "10001011", 8093 => "11111111", 8094 => "01000010", 8095 => "00110100", 8096 => "10001100", 8097 => "01100101", 8099 => "00101001", 8100 => "01000000", 8101 => "10011100", 8102 => "11101011", 8104 => "01111100", 8108 => "10010010", 8112 => "00111001", 8113 => "10100110", 8115 => "10010010", 8120 => "11101010", 8124 => "01101111", 8125 => "11000111", 8127 => "00101010", 8131 => "11100001", 8133 => "11111001", 8134 => "11111110", 8136 => "11101100", 8139 => "10111010", 8140 => "01100011", 8142 => "00010111", 8145 => "11011011", 8146 => "10001000", 8147 => "00110010", 8148 => "10000010", 8150 => "11111110", 8151 => "00001100", 8152 => "11001100", 8155 => "01101110", 8156 => "01111001", 8157 => "01000110", 8164 => "00011001", 8165 => "00000001", 8167 => "01010000", 8168 => "10000100", 8169 => "11111101", 8170 => "01011110", 8171 => "00000001", 8172 => "01100001", 8174 => "10010010", 8175 => "11011110", 8176 => "00110010", 8178 => "11101111", 8183 => "10110111", 8185 => "00010001", 8186 => "10001001", 8187 => "11010000", 8191 => "01111000", 8197 => "01001111", 8200 => "11000110", 8201 => "10011011", 8203 => "11101101", 8204 => "00111011", 8205 => "11001010", 8207 => "01011110", 8210 => "10101011", 8213 => "10100001", 8217 => "00011101", 8219 => "00101010", 8223 => "11011110", 8228 => "00111110", 8229 => "00001010", 8233 => "00010110", 8235 => "01111000", 8239 => "11000100", 8241 => "01111111", 8242 => "10110110", 8244 => "00111010", 8245 => "10010101", 8247 => "10101000", 8248 => "10000011", 8249 => "11111100", 8253 => "11111000", 8254 => "01100000", 8255 => "00100101", 8256 => "11001001", 8257 => "00010000", 8261 => "11110111", 8262 => "00100000", 8263 => "01110100", 8264 => "10011111", 8265 => "01011010", 8268 => "11110100", 8275 => "00110000", 8277 => "01010101", 8279 => "00111100", 8280 => "00111010", 8282 => "00101111", 8285 => "00010000", 8289 => "11110110", 8292 => "10001010", 8296 => "11110000", 8297 => "11001001", 8299 => "11000110", 8301 => "11001000", 8302 => "00101011", 8304 => "01011100", 8306 => "01010111", 8307 => "01111001", 8308 => "00000111", 8312 => "11110111", 8313 => "11101011", 8314 => "01011001", 8318 => "11100001", 8320 => "00000001", 8321 => "00100101", 8323 => "11000010", 8325 => "00101010", 8326 => "10110010", 8327 => "01010100", 8328 => "00110111", 8330 => "10110111", 8331 => "01010010", 8334 => "00101000", 8337 => "01101101", 8338 => "10110110", 8339 => "10001111", 8340 => "01010001", 8341 => "01111110", 8342 => "01101111", 8343 => "01111110", 8344 => "10001110", 8346 => "01110010", 8351 => "00010111", 8354 => "11001000", 8358 => "01010100", 8362 => "01000001", 8364 => "10001110", 8366 => "00101110", 8367 => "10000111", 8370 => "10001011", 8372 => "10010101", 8373 => "01010011", 8377 => "10101001", 8378 => "10100101", 8379 => "11110000", 8380 => "00001001", 8382 => "00000011", 8383 => "10110100", 8384 => "00111011", 8385 => "00001010", 8386 => "00011000", 8388 => "11000110", 8389 => "10100110", 8390 => "10011000", 8391 => "10010011", 8393 => "00101110", 8394 => "10110000", 8396 => "00011100", 8398 => "01011101", 8400 => "00100111", 8402 => "00110011", 8407 => "10011000", 8409 => "10011100", 8411 => "11100111", 8413 => "11100101", 8416 => "10000011", 8417 => "01111011", 8418 => "01000111", 8419 => "01101011", 8421 => "01111010", 8422 => "00111000", 8423 => "10101011", 8424 => "01101111", 8427 => "11010011", 8428 => "01101011", 8430 => "10100110", 8431 => "11100111", 8435 => "00101000", 8438 => "11101010", 8440 => "01010011", 8441 => "01110100", 8442 => "10101000", 8445 => "10010111", 8446 => "11000010", 8452 => "00101001", 8455 => "10110010", 8456 => "11110111", 8460 => "00001111", 8462 => "01100000", 8464 => "10011100", 8465 => "11011111", 8470 => "11001101", 8471 => "01101010", 8473 => "00110100", 8475 => "10111100", 8476 => "01010000", 8477 => "10011001", 8478 => "00001000", 8479 => "00111111", 8480 => "00100001", 8481 => "10011000", 8483 => "10010101", 8484 => "11100101", 8485 => "11111011", 8493 => "10010100", 8494 => "00011001", 8498 => "11110111", 8499 => "10000011", 8500 => "00101100", 8502 => "01110011", 8505 => "01011001", 8506 => "01100011", 8507 => "01000000", 8508 => "01001010", 8511 => "10011000", 8513 => "00111100", 8514 => "10010011", 8515 => "10010111", 8523 => "11110011", 8524 => "11110000", 8525 => "01000101", 8526 => "11011000", 8527 => "10101000", 8530 => "00101110", 8531 => "11110011", 8532 => "10111111", 8533 => "10001010", 8535 => "00100011", 8537 => "00010100", 8538 => "00000010", 8541 => "11010010", 8542 => "11010001", 8543 => "11010000", 8546 => "11000101", 8547 => "10011011", 8552 => "01110100", 8553 => "11011011", 8555 => "10010001", 8560 => "01110100", 8561 => "01110001", 8562 => "01110101", 8563 => "10010010", 8565 => "10110010", 8566 => "11111100", 8567 => "00111011", 8568 => "11100000", 8570 => "11001100", 8571 => "10001100", 8572 => "11000100", 8574 => "10100110", 8576 => "11001101", 8577 => "10100101", 8578 => "10001001", 8585 => "01101000", 8586 => "10000100", 8587 => "00010001", 8591 => "01001001", 8595 => "01011100", 8596 => "01110100", 8598 => "10010110", 8599 => "10010100", 8600 => "11001001", 8602 => "00101011", 8603 => "00010000", 8604 => "00001010", 8607 => "10111011", 8609 => "11111010", 8612 => "10011011", 8613 => "10111000", 8614 => "01001111", 8615 => "01100000", 8616 => "10000110", 8617 => "01001101", 8620 => "11011000", 8621 => "00001101", 8622 => "00110111", 8625 => "00000101", 8628 => "11011011", 8633 => "11011111", 8641 => "11010110", 8645 => "11111010", 8648 => "01100011", 8651 => "01001010", 8655 => "00101010", 8656 => "00010001", 8658 => "00101100", 8662 => "00001001", 8664 => "00110101", 8667 => "10010010", 8669 => "10001100", 8670 => "01001000", 8672 => "00000010", 8673 => "00000001", 8674 => "11010100", 8676 => "00000010", 8677 => "01001110", 8680 => "01110101", 8681 => "00111100", 8683 => "11011011", 8685 => "11101101", 8689 => "00000111", 8691 => "01011010", 8693 => "01110010", 8694 => "10110101", 8695 => "00000111", 8698 => "10010011", 8700 => "00001001", 8701 => "10110010", 8703 => "10100010", 8705 => "10111101", 8706 => "00110010", 8707 => "10100100", 8710 => "11000000", 8713 => "00001100", 8715 => "10101010", 8717 => "11111001", 8721 => "10110001", 8723 => "11100110", 8725 => "00000001", 8727 => "01001110", 8728 => "10010011", 8729 => "01011000", 8731 => "10000011", 8734 => "01011011", 8737 => "10010101", 8738 => "00010000", 8739 => "11110110", 8740 => "01110001", 8742 => "10001001", 8747 => "11001101", 8748 => "01011000", 8751 => "01111010", 8752 => "01001010", 8755 => "01110100", 8758 => "11101101", 8762 => "00010001", 8763 => "01011110", 8765 => "11101101", 8768 => "00111001", 8770 => "01110100", 8771 => "01001101", 8773 => "01110100", 8774 => "00101100", 8775 => "00001100", 8776 => "00011010", 8777 => "00011101", 8779 => "10111001", 8783 => "10110110", 8784 => "11111000", 8787 => "00110111", 8796 => "11011011", 8798 => "00100111", 8801 => "01011100", 8803 => "00001011", 8804 => "01011111", 8809 => "10110100", 8813 => "01100111", 8817 => "11111001", 8822 => "00110000", 8825 => "11100000", 8826 => "10111101", 8827 => "01010111", 8831 => "00000100", 8832 => "10000111", 8833 => "11001000", 8834 => "10110111", 8836 => "01101110", 8839 => "01111010", 8840 => "10000101", 8844 => "10000001", 8846 => "01010100", 8847 => "00110001", 8848 => "10010100", 8852 => "10111000", 8854 => "11110000", 8856 => "01100101", 8857 => "10110000", 8859 => "00001100", 8860 => "10110110", 8861 => "10011100", 8863 => "11011110", 8864 => "10100110", 8867 => "00001001", 8869 => "01111011", 8870 => "00111101", 8871 => "10001010", 8873 => "00000110", 8876 => "00111001", 8877 => "01110101", 8878 => "11110001", 8880 => "10101010", 8881 => "00100110", 8882 => "11000001", 8883 => "10110000", 8885 => "01000001", 8887 => "11101010", 8888 => "11000100", 8889 => "01101010", 8890 => "00110110", 8893 => "01011110", 8894 => "01101011", 8895 => "01111000", 8897 => "01001100", 8898 => "10111001", 8904 => "10111011", 8916 => "01100001", 8917 => "01000011", 8921 => "10010010", 8927 => "00011000", 8931 => "01001111", 8932 => "00101010", 8933 => "00100001", 8938 => "01100101", 8939 => "00110110", 8940 => "10101000", 8941 => "01100110", 8945 => "01100111", 8951 => "00000111", 8952 => "11100010", 8954 => "10000011", 8955 => "11100101", 8956 => "11111011", 8957 => "10100010", 8959 => "10111100", 8960 => "00000110", 8962 => "00011011", 8966 => "01011001", 8967 => "00111010", 8971 => "11000111", 8976 => "11101101", 8977 => "01101011", 8979 => "10010101", 8980 => "00000111", 8982 => "10000101", 8988 => "01100000", 8989 => "10010011", 8991 => "10011011", 8992 => "11100000", 8994 => "00111001", 9007 => "10110110", 9009 => "00110111", 9010 => "10000001", 9011 => "11100011", 9013 => "01111001", 9014 => "10111101", 9015 => "10011011", 9017 => "10100101", 9018 => "00100011", 9019 => "00111010", 9023 => "10010011", 9030 => "11000111", 9035 => "11110001", 9036 => "10111111", 9037 => "00001101", 9038 => "11011000", 9039 => "10011000", 9040 => "01111111", 9042 => "10100010", 9044 => "00001100", 9045 => "01000110", 9049 => "10101100", 9050 => "00011000", 9052 => "00001100", 9057 => "00111001", 9061 => "11111100", 9063 => "00010000", 9064 => "11111110", 9065 => "11011011", 9066 => "10101001", 9067 => "01100101", 9068 => "00100011", 9071 => "01111101", 9072 => "11101100", 9073 => "00100100", 9074 => "00110001", 9075 => "00111101", 9076 => "01101000", 9082 => "11000101", 9083 => "00011010", 9084 => "11011100", 9085 => "11010100", 9086 => "00001111", 9089 => "01101001", 9092 => "01100010", 9093 => "10111111", 9096 => "01101000", 9101 => "11010101", 9102 => "01101000", 9105 => "10111011", 9107 => "00100010", 9109 => "11111010", 9110 => "01111001", 9111 => "00101110", 9112 => "01010101", 9115 => "00001010", 9116 => "00100100", 9117 => "10100111", 9119 => "01101010", 9120 => "10110010", 9121 => "01101000", 9123 => "01110101", 9125 => "11100011", 9127 => "11101111", 9129 => "00101011", 9133 => "01011010", 9135 => "01010001", 9137 => "10100000", 9144 => "01010100", 9145 => "10100000", 9146 => "10010111", 9147 => "01110110", 9150 => "01011110", 9152 => "00101100", 9153 => "00001110", 9154 => "10010101", 9155 => "11111011", 9156 => "10101111", 9157 => "11110101", 9158 => "00001111", 9159 => "11100110", 9162 => "10010010", 9163 => "01010101", 9166 => "11000100", 9169 => "11000000", 9173 => "10111101", 9174 => "10111001", 9176 => "10100111", 9179 => "10110110", 9181 => "10011011", 9185 => "00110100", 9187 => "10000111", 9192 => "10110101", 9195 => "00010100", 9196 => "11101010", 9198 => "11011110", 9199 => "10111001", 9202 => "01111001", 9203 => "11001110", 9204 => "01011010", 9205 => "01101100", 9206 => "11110110", 9208 => "01001111", 9211 => "10110001", 9212 => "01000110", 9214 => "10001100", 9215 => "10010000", 9216 => "00000101", 9217 => "11111011", 9220 => "01100111", 9221 => "01001110", 9222 => "01010101", 9223 => "11110111", 9226 => "01000111", 9230 => "00100100", 9232 => "00000100", 9233 => "01001100", 9238 => "01001101", 9239 => "00001001", 9240 => "00101110", 9242 => "01000110", 9247 => "10010001", 9249 => "00010010", 9252 => "10111010", 9253 => "11101110", 9255 => "01000000", 9256 => "10110100", 9257 => "01010110", 9258 => "11101010", 9259 => "01011101", 9263 => "11101000", 9265 => "01010001", 9267 => "10100111", 9268 => "01001001", 9269 => "10101010", 9270 => "00010111", 9271 => "11101011", 9274 => "01101000", 9278 => "10010111", 9279 => "00001011", 9280 => "10010000", 9283 => "01111001", 9284 => "11000001", 9285 => "01011001", 9286 => "10000010", 9288 => "01000011", 9290 => "11101010", 9293 => "10010001", 9294 => "00010011", 9295 => "00010101", 9297 => "10100111", 9298 => "01110100", 9299 => "01110111", 9301 => "11101101", 9303 => "10101001", 9305 => "01001000", 9306 => "01100011", 9307 => "10001100", 9309 => "00101010", 9312 => "10001010", 9313 => "10011001", 9315 => "01000100", 9317 => "10001000", 9320 => "01101010", 9321 => "11010110", 9323 => "00110000", 9324 => "01100100", 9325 => "10111110", 9326 => "01010111", 9329 => "00101011", 9330 => "11110000", 9331 => "10010111", 9333 => "01110100", 9336 => "00011110", 9337 => "11000011", 9342 => "01001010", 9343 => "01001010", 9344 => "11011110", 9345 => "10110110", 9348 => "11110100", 9349 => "00011100", 9350 => "10111011", 9352 => "10010001", 9353 => "10010000", 9357 => "00011111", 9366 => "00110001", 9368 => "11111010", 9369 => "00011100", 9370 => "11100001", 9371 => "00100100", 9373 => "00000010", 9376 => "00111100", 9377 => "00000101", 9379 => "11100100", 9380 => "11110101", 9384 => "11000011", 9386 => "00001010", 9387 => "01110111", 9390 => "10110111", 9391 => "00010111", 9392 => "01111111", 9393 => "00011111", 9395 => "10111100", 9396 => "11111001", 9397 => "00001011", 9398 => "01010000", 9404 => "00011001", 9406 => "00101101", 9408 => "10101011", 9410 => "10010111", 9418 => "11110111", 9420 => "11110000", 9422 => "10101000", 9424 => "01110001", 9429 => "01011110", 9435 => "01111001", 9437 => "00101001", 9438 => "10001101", 9439 => "00101011", 9440 => "11001101", 9443 => "11110011", 9447 => "11101100", 9450 => "11010110", 9453 => "11011100", 9454 => "11111001", 9456 => "11000000", 9457 => "01011001", 9460 => "10111110", 9461 => "01100101", 9463 => "11000011", 9464 => "00011111", 9466 => "01010010", 9467 => "10010000", 9469 => "11000110", 9470 => "01101101", 9474 => "01001111", 9477 => "01101111", 9478 => "11011101", 9480 => "00100100", 9481 => "10001001", 9484 => "10100101", 9486 => "00111110", 9488 => "10011100", 9490 => "11111010", 9491 => "01111101", 9494 => "01100000", 9497 => "11000010", 9500 => "11111001", 9502 => "00100101", 9504 => "10000111", 9505 => "00011101", 9507 => "01110110", 9510 => "01000000", 9511 => "00010110", 9513 => "00110100", 9516 => "10011010", 9518 => "01000110", 9519 => "11010000", 9520 => "11110101", 9522 => "10001101", 9524 => "01000010", 9525 => "00111011", 9526 => "01101000", 9527 => "00100010", 9529 => "11100100", 9530 => "10001111", 9532 => "00111011", 9533 => "11001100", 9534 => "11011010", 9537 => "10101001", 9545 => "00000101", 9547 => "10000101", 9549 => "01111010", 9550 => "01111110", 9552 => "10010110", 9553 => "01010011", 9554 => "00110100", 9555 => "10100010", 9556 => "10010110", 9557 => "01110011", 9558 => "00101111", 9559 => "10000011", 9560 => "11111011", 9562 => "01001100", 9564 => "00100000", 9565 => "10101100", 9568 => "10000010", 9569 => "00101111", 9571 => "11111111", 9572 => "10110101", 9575 => "01000101", 9578 => "01111010", 9579 => "11011110", 9580 => "01110001", 9583 => "00001010", 9584 => "01111111", 9587 => "00001000", 9592 => "11101000", 9601 => "00101110", 9602 => "11011110", 9603 => "01010010", 9604 => "00001001", 9606 => "01110110", 9607 => "01010101", 9609 => "01111101", 9610 => "01010110", 9611 => "01101010", 9616 => "10001101", 9619 => "00100110", 9621 => "11001000", 9623 => "00001010", 9624 => "01100111", 9626 => "10011011", 9628 => "11100100", 9629 => "00011101", 9630 => "10110010", 9632 => "11111100", 9634 => "11101000", 9639 => "01100000", 9640 => "01000011", 9642 => "11011000", 9647 => "11110001", 9651 => "00101111", 9656 => "01010111", 9660 => "10110000", 9661 => "01100110", 9662 => "11011111", 9663 => "11011101", 9665 => "10010001", 9671 => "10011110", 9675 => "11000010", 9676 => "00110001", 9678 => "11010100", 9679 => "01111110", 9681 => "10010011", 9683 => "00101100", 9685 => "01111101", 9686 => "10111000", 9688 => "01111011", 9689 => "00001000", 9691 => "00100000", 9693 => "11010011", 9696 => "11111011", 9701 => "10101011", 9702 => "00010011", 9706 => "01110000", 9710 => "10110011", 9711 => "10011011", 9712 => "00111001", 9716 => "10111001", 9719 => "11001001", 9720 => "11001100", 9722 => "00001001", 9725 => "01111101", 9730 => "01001001", 9733 => "00110110", 9734 => "01011001", 9739 => "00101000", 9742 => "10001111", 9746 => "11010001", 9748 => "01110000", 9751 => "01001000", 9752 => "11011100", 9753 => "00100010", 9757 => "10000000", 9758 => "10000000", 9762 => "01110000", 9763 => "11101001", 9765 => "01000010", 9771 => "11010111", 9773 => "00000001", 9777 => "10011001", 9780 => "11011011", 9781 => "10001101", 9783 => "10011000", 9784 => "01111000", 9786 => "11111001", 9789 => "10111011", 9790 => "00011111", 9791 => "10111001", 9794 => "11110101", 9796 => "00100101", 9797 => "01001111", 9798 => "10010101", 9803 => "01111001", 9804 => "10001110", 9806 => "00100001", 9807 => "01100011", 9808 => "01011010", 9809 => "11111101", 9811 => "11000011", 9814 => "11110111", 9819 => "10111011", 9820 => "11000111", 9824 => "01011010", 9825 => "00101011", 9826 => "00011111", 9833 => "10000001", 9834 => "00010111", 9836 => "00011100", 9837 => "10000000", 9842 => "01110100", 9843 => "00111000", 9845 => "10100110", 9847 => "00011010", 9848 => "00110001", 9851 => "00101011", 9852 => "01111110", 9853 => "00111011", 9854 => "01011100", 9856 => "11001001", 9857 => "00001110", 9858 => "10111011", 9859 => "11010110", 9860 => "01101100", 9863 => "10100001", 9866 => "00100100", 9867 => "11100100", 9868 => "00100110", 9873 => "01011110", 9876 => "01010101", 9878 => "01011111", 9881 => "00100110", 9882 => "11110110", 9884 => "01000000", 9885 => "10000011", 9891 => "10000001", 9892 => "01110101", 9893 => "00111110", 9897 => "01100001", 9898 => "10111001", 9900 => "01110011", 9902 => "00010110", 9903 => "00001100", 9911 => "10000011", 9912 => "01101010", 9913 => "01000101", 9917 => "10110010", 9918 => "11011100", 9921 => "00110101", 9922 => "01011101", 9923 => "11000000", 9925 => "00111110", 9927 => "01110110", 9928 => "01011001", 9930 => "10100011", 9931 => "00011101", 9932 => "10001111", 9933 => "10111101", 9938 => "11111101", 9946 => "11111100", 9947 => "00110001", 9950 => "00011000", 9962 => "10110010", 9963 => "10110001", 9965 => "01100110", 9967 => "00101101", 9970 => "00110011", 9973 => "01001110", 9975 => "00110100", 9976 => "11111001", 9978 => "11000101", 9982 => "10011100", 9983 => "00001101", 9986 => "11111111", 9988 => "11010010", 9989 => "00011010", 9990 => "10100101", 9992 => "11000100", 9995 => "01101000", 9996 => "00010001", 9999 => "00101011", 10000 => "11011011", 10001 => "00000010", 10002 => "10010010", 10005 => "10110001", 10008 => "00011001", 10014 => "11101100", 10016 => "11010001", 10018 => "11110011", 10025 => "10011010", 10026 => "10010011", 10030 => "11000000", 10033 => "11001011", 10034 => "00100010", 10038 => "10001010", 10039 => "01101110", 10043 => "10000000", 10044 => "00011111", 10045 => "10100001", 10046 => "01110000", 10047 => "11000110", 10048 => "01110000", 10050 => "00001110", 10052 => "01101101", 10055 => "11000011", 10056 => "11111100", 10057 => "00101001", 10059 => "10100000", 10062 => "11111000", 10063 => "00101111", 10064 => "00101011", 10066 => "10010110", 10067 => "11000111", 10070 => "00010000", 10078 => "00101010", 10079 => "00100011", 10086 => "10000111", 10090 => "11101011", 10091 => "00110111", 10093 => "01001110", 10096 => "11001110", 10098 => "11111001", 10099 => "11010000", 10101 => "10111010", 10102 => "10111101", 10103 => "01000000", 10105 => "11111100", 10107 => "10110111", 10108 => "00100001", 10109 => "00111110", 10110 => "11000010", 10111 => "00110101", 10113 => "01110100", 10117 => "11010011", 10119 => "01100010", 10120 => "10101010", 10125 => "10100111", 10127 => "10111001", 10128 => "01010011", 10129 => "00010011", 10131 => "00101110", 10133 => "00001100", 10134 => "10100001", 10136 => "00011110", 10137 => "10010000", 10141 => "00111110", 10142 => "10101000", 10144 => "11010000", 10147 => "00101110", 10149 => "00101100", 10150 => "10000011", 10154 => "00110000", 10157 => "10000011", 10158 => "10111110", 10159 => "10100110", 10160 => "10110111", 10162 => "01100011", 10165 => "01011000", 10166 => "11110001", 10168 => "11010000", 10169 => "01000110", 10170 => "01000010", 10172 => "01110100", 10173 => "11101111", 10176 => "10101001", 10178 => "00010010", 10180 => "10001100", 10181 => "10001111", 10182 => "00011110", 10184 => "11110001", 10185 => "10100000", 10186 => "00101101", 10188 => "00110111", 10189 => "10110011", 10191 => "01110001", 10196 => "11100100", 10198 => "00110110", 10199 => "10011001", 10201 => "00011010", 10202 => "00100111", 10206 => "11101000", 10209 => "00101011", 10210 => "11011001", 10211 => "11011100", 10219 => "00010111", 10222 => "01101101", 10229 => "00101100", 10231 => "11000111", 10233 => "01001001", 10235 => "01100110", 10236 => "10111010", 10238 => "00101000", 10240 => "00110100", 10242 => "11010100", 10243 => "10011111", 10246 => "00111110", 10248 => "01101011", 10250 => "11000110", 10251 => "10011110", 10252 => "00101011", 10253 => "00100111", 10254 => "01001101", 10255 => "10010010", 10257 => "11101010", 10259 => "11010001", 10262 => "01010000", 10263 => "11000111", 10265 => "00001100", 10268 => "11111001", 10270 => "11101111", 10271 => "01111001", 10274 => "00000001", 10276 => "01011111", 10280 => "01110000", 10284 => "00001100", 10287 => "01100111", 10288 => "01110001", 10290 => "10000001", 10291 => "10110111", 10293 => "11011110", 10295 => "01101101", 10296 => "11001001", 10297 => "01011110", 10300 => "00110110", 10301 => "01001110", 10303 => "10011111", 10304 => "11000100", 10306 => "01101110", 10307 => "01000001", 10308 => "10111011", 10310 => "10111000", 10311 => "10001100", 10313 => "01001000", 10314 => "01110011", 10315 => "10111010", 10319 => "11110111", 10321 => "11110110", 10322 => "10100101", 10323 => "00000001", 10324 => "10001110", 10327 => "10010110", 10331 => "01001111", 10332 => "01000001", 10333 => "00110101", 10334 => "10100001", 10336 => "11101001", 10337 => "11111001", 10342 => "10011011", 10345 => "01101111", 10347 => "11001001", 10350 => "10000000", 10352 => "10000110", 10353 => "11101110", 10355 => "11111010", 10356 => "01111010", 10359 => "10110110", 10362 => "11011111", 10364 => "10110110", 10365 => "00111101", 10366 => "00010011", 10369 => "00110000", 10370 => "11010011", 10371 => "01111100", 10374 => "11101000", 10375 => "10011010", 10377 => "10100000", 10378 => "00011010", 10381 => "10001000", 10382 => "11100111", 10389 => "00011100", 10395 => "11011001", 10396 => "01100111", 10397 => "01000110", 10401 => "10001100", 10402 => "11010001", 10407 => "10000101", 10409 => "01100010", 10412 => "10100111", 10414 => "10111001", 10415 => "00110010", 10416 => "01011111", 10417 => "10000001", 10419 => "01011111", 10421 => "11001100", 10422 => "11000001", 10423 => "00100010", 10424 => "10101001", 10426 => "10001010", 10427 => "10010000", 10430 => "11100111", 10431 => "11100110", 10432 => "10010111", 10433 => "10100011", 10435 => "01000011", 10436 => "01011101", 10439 => "01010111", 10443 => "01010111", 10447 => "10100000", 10454 => "00000101", 10456 => "10101011", 10458 => "10100011", 10461 => "11000110", 10462 => "10011100", 10464 => "11111101", 10466 => "10000000", 10468 => "01010010", 10469 => "00001000", 10472 => "00100010", 10475 => "01010000", 10479 => "01001100", 10480 => "11111110", 10482 => "11101111", 10483 => "00001100", 10486 => "00101101", 10487 => "10101001", 10490 => "10010001", 10492 => "00100001", 10493 => "01011100", 10495 => "01110010", 10501 => "11101011", 10502 => "11101011", 10503 => "00000111", 10505 => "01110101", 10506 => "10011110", 10507 => "00011101", 10508 => "10001100", 10509 => "10011000", 10510 => "11000100", 10511 => "01100000", 10512 => "10001010", 10517 => "00110000", 10520 => "10010111", 10521 => "00110111", 10524 => "00111010", 10526 => "01110111", 10527 => "00001000", 10528 => "10110000", 10530 => "10000100", 10531 => "01001010", 10532 => "11100010", 10533 => "01110010", 10534 => "00000110", 10537 => "11111000", 10539 => "01010010", 10541 => "11011001", 10542 => "00011000", 10544 => "01101010", 10545 => "11000010", 10548 => "00100111", 10552 => "11000010", 10553 => "10100011", 10555 => "00101100", 10557 => "10011010", 10558 => "01001010", 10559 => "11000101", 10561 => "11000110", 10562 => "01000001", 10564 => "00111001", 10565 => "11010001", 10567 => "11111011", 10570 => "11011001", 10572 => "10000000", 10573 => "11010001", 10575 => "10011011", 10577 => "00101000", 10579 => "01001000", 10581 => "10010010", 10583 => "01101111", 10584 => "01110101", 10585 => "11011000", 10586 => "00011010", 10587 => "00110000", 10589 => "10110001", 10590 => "01001110", 10594 => "11000000", 10596 => "01011001", 10598 => "00011101", 10601 => "00101010", 10602 => "01100111", 10604 => "10101000", 10608 => "11001011", 10610 => "10001111", 10612 => "01010110", 10613 => "01111111", 10614 => "10110001", 10615 => "00111101", 10618 => "10100100", 10619 => "01001010", 10620 => "01011000", 10621 => "00000011", 10622 => "00110101", 10624 => "00110000", 10626 => "10010011", 10627 => "11000011", 10628 => "00011100", 10630 => "11101010", 10631 => "00001010", 10632 => "11110011", 10633 => "10101101", 10636 => "11000011", 10637 => "01111001", 10638 => "11011010", 10639 => "00100110", 10640 => "01110011", 10641 => "01010000", 10647 => "11100001", 10648 => "11100000", 10650 => "00110110", 10651 => "11001111", 10652 => "00101111", 10653 => "10110000", 10654 => "00000010", 10656 => "01011100", 10657 => "10110110", 10658 => "11101001", 10660 => "10010101", 10663 => "01011110", 10664 => "11010101", 10667 => "01000000", 10668 => "11010011", 10672 => "10011110", 10674 => "10001100", 10675 => "11110000", 10677 => "01000111", 10679 => "11011011", 10680 => "00100111", 10681 => "11010010", 10683 => "00101010", 10684 => "00010111", 10686 => "11101001", 10687 => "11001101", 10693 => "01001110", 10698 => "11111101", 10700 => "01101100", 10701 => "01000100", 10704 => "01010001", 10706 => "01001000", 10708 => "11111001", 10709 => "11011111", 10710 => "00000011", 10713 => "10001011", 10716 => "10000010", 10722 => "11110101", 10723 => "10110010", 10724 => "11011011", 10725 => "11100000", 10727 => "01010101", 10733 => "00011000", 10734 => "00000100", 10735 => "11010110", 10739 => "11000010", 10741 => "00101100", 10742 => "00110110", 10744 => "11011100", 10745 => "01100111", 10746 => "10110111", 10748 => "10100001", 10750 => "11010010", 10752 => "10101011", 10753 => "10000100", 10754 => "01100001", 10755 => "00100010", 10760 => "01000101", 10765 => "01010100", 10766 => "01000110", 10767 => "00011110", 10768 => "01110000", 10769 => "11000101", 10772 => "00001110", 10774 => "01111001", 10775 => "00010111", 10777 => "11000100", 10779 => "01011100", 10783 => "01011111", 10784 => "01001010", 10785 => "00111001", 10786 => "00011001", 10793 => "01010100", 10794 => "00100011", 10795 => "01100000", 10798 => "11101100", 10799 => "11000100", 10801 => "01101101", 10808 => "00011110", 10811 => "11110100", 10815 => "11100100", 10816 => "10100010", 10818 => "11110001", 10819 => "11110101", 10821 => "11010010", 10823 => "01110011", 10826 => "00001110", 10828 => "01001011", 10829 => "00010011", 10831 => "10110100", 10834 => "01101100", 10835 => "11101010", 10836 => "01001000", 10838 => "00010101", 10839 => "10001111", 10841 => "00000111", 10843 => "01000011", 10844 => "11011001", 10847 => "01110001", 10849 => "00101100", 10850 => "10000011", 10852 => "01110011", 10853 => "11111101", 10854 => "11110011", 10855 => "01001110", 10857 => "11101010", 10861 => "10101010", 10862 => "01110010", 10863 => "10110000", 10867 => "10001110", 10868 => "01000000", 10869 => "10100111", 10871 => "11011010", 10872 => "00100010", 10874 => "11100101", 10875 => "00100101", 10876 => "10001010", 10877 => "00000010", 10881 => "00000101", 10882 => "00110010", 10883 => "10010010", 10885 => "10010001", 10886 => "10011000", 10887 => "00110101", 10888 => "11010000", 10889 => "11111101", 10890 => "10100111", 10893 => "10000111", 10895 => "11001101", 10896 => "00000100", 10897 => "01010101", 10898 => "00101100", 10902 => "10101100", 10903 => "00001110", 10905 => "11101000", 10907 => "01010000", 10908 => "11010100", 10917 => "00001000", 10919 => "00100001", 10920 => "10111101", 10923 => "11001101", 10924 => "01001000", 10926 => "11110000", 10928 => "01011100", 10931 => "10110010", 10936 => "00000111", 10937 => "11010100", 10938 => "00010001", 10939 => "11011111", 10941 => "11010010", 10943 => "11011000", 10944 => "11000101", 10945 => "10011010", 10946 => "01110110", 10949 => "11000010", 10950 => "10000100", 10954 => "01001111", 10955 => "11111011", 10956 => "00101000", 10957 => "01011110", 10959 => "00001001", 10963 => "10010101", 10966 => "10011010", 10967 => "00100010", 10968 => "11100110", 10969 => "01010111", 10972 => "00110111", 10973 => "11101100", 10976 => "00100000", 10978 => "00010100", 10979 => "10010110", 10980 => "00100001", 10983 => "01011100", 10984 => "11100011", 10985 => "11101011", 10986 => "10000111", 10988 => "11010110", 10990 => "10101000", 10994 => "00010110", 10996 => "01010101", 11001 => "00110010", 11003 => "10011111", 11004 => "01011110", 11005 => "00101111", 11006 => "10011111", 11009 => "01000111", 11012 => "01110110", 11014 => "11100111", 11016 => "11000110", 11025 => "10011111", 11026 => "10101101", 11027 => "11110011", 11028 => "10000010", 11031 => "10010010", 11034 => "11011101", 11035 => "11011000", 11038 => "00000100", 11045 => "01010101", 11046 => "10010000", 11048 => "11011100", 11049 => "00000111", 11051 => "00101010", 11052 => "11101001", 11053 => "10101100", 11054 => "01110111", 11055 => "10010001", 11056 => "01110110", 11059 => "11011111", 11060 => "00010101", 11061 => "00110111", 11065 => "01101011", 11069 => "01100010", 11071 => "01001010", 11072 => "00000100", 11073 => "00000010", 11074 => "11111000", 11075 => "00011101", 11076 => "11100100", 11077 => "01101010", 11078 => "00010111", 11079 => "11111011", 11080 => "10010101", 11081 => "11110110", 11082 => "10000100", 11084 => "10101110", 11087 => "00101100", 11088 => "11011110", 11090 => "00100010", 11093 => "01000101", 11094 => "11011010", 11096 => "11001110", 11099 => "10111111", 11103 => "01001011", 11106 => "01110001", 11107 => "11100101", 11111 => "11100000", 11113 => "00101101", 11114 => "10110010", 11115 => "01011100", 11119 => "11101000", 11120 => "11011011", 11125 => "10001100", 11126 => "01110011", 11127 => "10011011", 11128 => "01010011", 11130 => "10101011", 11133 => "10111101", 11134 => "00100101", 11136 => "00010010", 11137 => "01110101", 11138 => "10011101", 11139 => "00010100", 11141 => "00100001", 11142 => "01111000", 11143 => "00111000", 11145 => "11001101", 11148 => "10101101", 11150 => "01101010", 11151 => "10111000", 11154 => "11000110", 11158 => "00111101", 11160 => "01110100", 11162 => "00110110", 11164 => "00001111", 11165 => "00010001", 11170 => "10110011", 11177 => "10110101", 11178 => "00100000", 11181 => "01010010", 11183 => "00111010", 11184 => "11011011", 11187 => "01100010", 11190 => "10100000", 11192 => "10101011", 11195 => "11010111", 11196 => "01001011", 11199 => "00110110", 11203 => "01011001", 11206 => "01001011", 11210 => "00000010", 11213 => "11110111", 11219 => "00000001", 11220 => "00010001", 11221 => "11111001", 11222 => "00111101", 11226 => "11100010", 11229 => "00010010", 11232 => "00000010", 11233 => "10001100", 11237 => "10110111", 11238 => "10111011", 11239 => "11111101", 11241 => "10010100", 11242 => "10000101", 11243 => "10110000", 11248 => "11010101", 11249 => "11001100", 11250 => "00111011", 11252 => "01101110", 11254 => "00011100", 11255 => "01011011", 11257 => "00000100", 11258 => "11101010", 11259 => "11110010", 11261 => "00000001", 11264 => "01101101", 11265 => "11110011", 11266 => "11100111", 11267 => "00101000", 11270 => "00001011", 11271 => "10010111", 11273 => "10000110", 11274 => "10011111", 11275 => "10010101", 11276 => "01100111", 11277 => "01000010", 11279 => "00011101", 11280 => "01001010", 11281 => "11011011", 11284 => "10011001", 11285 => "10011100", 11286 => "11000000", 11288 => "01101111", 11293 => "00011001", 11296 => "10101001", 11297 => "00011000", 11298 => "01000000", 11300 => "00010101", 11301 => "10001011", 11302 => "01101000", 11303 => "10101100", 11304 => "00100111", 11306 => "01101111", 11307 => "11000101", 11309 => "00111010", 11311 => "10111011", 11312 => "00110011", 11313 => "00101111", 11316 => "00000100", 11318 => "11011001", 11320 => "01010000", 11322 => "00000011", 11323 => "10010111", 11326 => "10001001", 11327 => "11101111", 11329 => "10000001", 11330 => "11100101", 11336 => "01111110", 11337 => "01000110", 11339 => "11000100", 11342 => "11001000", 11343 => "11100111", 11345 => "01100111", 11347 => "10010110", 11348 => "00011001", 11349 => "01011011", 11350 => "00011001", 11351 => "00011111", 11352 => "01110010", 11353 => "01111011", 11358 => "00001101", 11363 => "10101010", 11365 => "10110111", 11366 => "10100000", 11367 => "11111011", 11368 => "10100100", 11369 => "10000111", 11371 => "11111100", 11373 => "10001100", 11374 => "01100010", 11376 => "10011001", 11377 => "00111101", 11378 => "11101001", 11382 => "11111010", 11385 => "01111111", 11386 => "01011110", 11387 => "11100101", 11388 => "11011100", 11391 => "01101101", 11392 => "01011101", 11394 => "01000000", 11395 => "11100010", 11396 => "01100110", 11398 => "11011100", 11400 => "00011011", 11404 => "01010100", 11407 => "00111001", 11408 => "01111011", 11409 => "11111100", 11411 => "10110100", 11413 => "01101000", 11415 => "01110001", 11416 => "11001000", 11417 => "01010011", 11422 => "10011111", 11423 => "01010101", 11424 => "10000001", 11425 => "01110101", 11426 => "00010110", 11429 => "01101110", 11431 => "11100100", 11432 => "11011110", 11434 => "11000101", 11435 => "11111110", 11437 => "10010111", 11438 => "00111100", 11440 => "11010110", 11441 => "01110011", 11442 => "01000111", 11443 => "01111000", 11444 => "11000101", 11445 => "10101100", 11447 => "11000110", 11448 => "10011101", 11449 => "10010011", 11450 => "01110000", 11451 => "11101110", 11453 => "00110111", 11454 => "01001110", 11455 => "11010011", 11457 => "11110100", 11458 => "11100011", 11460 => "00000011", 11461 => "10110001", 11469 => "00111111", 11479 => "01101010", 11480 => "10010000", 11483 => "11100010", 11486 => "10101000", 11487 => "10010010", 11488 => "11101110", 11489 => "01000000", 11490 => "10110110", 11492 => "01110011", 11494 => "01111101", 11495 => "01101100", 11499 => "01000001", 11502 => "01010000", 11504 => "10001110", 11506 => "00011011", 11507 => "10101001", 11508 => "00100111", 11511 => "00000100", 11513 => "10110010", 11517 => "01000101", 11519 => "10001100", 11520 => "11100101", 11522 => "11101011", 11524 => "11010110", 11528 => "11110010", 11532 => "10010101", 11534 => "11001100", 11537 => "00110010", 11540 => "00110111", 11541 => "01011010", 11545 => "00010000", 11547 => "11000111", 11548 => "10000101", 11549 => "00110011", 11550 => "11000111", 11552 => "10111000", 11553 => "11110110", 11554 => "10101001", 11555 => "01110011", 11557 => "01011001", 11562 => "11110100", 11564 => "00110100", 11565 => "01010011", 11567 => "00101010", 11568 => "00101001", 11569 => "10001111", 11572 => "11000000", 11573 => "11100110", 11574 => "11100001", 11576 => "10001000", 11577 => "11010000", 11578 => "10110010", 11579 => "11100011", 11585 => "01100100", 11587 => "00100101", 11588 => "11001111", 11592 => "10111011", 11596 => "11110110", 11601 => "11010101", 11602 => "01000010", 11604 => "01000001", 11605 => "10100000", 11606 => "01011001", 11607 => "01110011", 11611 => "10100001", 11612 => "00100101", 11613 => "10010101", 11618 => "00001100", 11620 => "00111010", 11622 => "00101111", 11623 => "00101000", 11624 => "10110100", 11625 => "11000001", 11627 => "00111110", 11628 => "01010101", 11632 => "01011110", 11634 => "10101010", 11635 => "10110110", 11637 => "11000010", 11639 => "10111000", 11640 => "01011001", 11641 => "10100100", 11643 => "10000000", 11652 => "11110110", 11656 => "10001100", 11659 => "01011001", 11664 => "11100001", 11665 => "10011110", 11667 => "11101110", 11668 => "00010010", 11669 => "00110001", 11671 => "01101101", 11672 => "00101000", 11673 => "11100011", 11674 => "00011100", 11675 => "01010010", 11676 => "01001100", 11679 => "01111000", 11681 => "00100110", 11683 => "11101111", 11684 => "10001101", 11687 => "11011100", 11691 => "10100010", 11693 => "00000111", 11700 => "01110100", 11701 => "00001000", 11703 => "00101110", 11704 => "11110110", 11706 => "01011001", 11707 => "01101101", 11708 => "10001101", 11709 => "00001001", 11710 => "00011000", 11711 => "00010110", 11712 => "00001100", 11713 => "00111111", 11715 => "11001011", 11717 => "01010011", 11720 => "10110100", 11723 => "00101100", 11724 => "01101010", 11725 => "11101111", 11726 => "10100101", 11727 => "00000011", 11728 => "00011111", 11735 => "11110000", 11737 => "00111010", 11742 => "00101010", 11745 => "01101111", 11746 => "11010010", 11747 => "01100110", 11748 => "11100100", 11749 => "11011110", 11752 => "01110100", 11753 => "11000001", 11755 => "11001011", 11760 => "10000101", 11761 => "01100000", 11762 => "01000100", 11764 => "11000000", 11766 => "01110000", 11767 => "10000101", 11769 => "00011110", 11770 => "00111011", 11771 => "10110111", 11773 => "10101011", 11776 => "11011011", 11778 => "11001011", 11779 => "00110111", 11781 => "01101000", 11782 => "01000001", 11783 => "11000101", 11784 => "11111010", 11785 => "01101001", 11787 => "01001110", 11791 => "10101101", 11792 => "10001111", 11793 => "10110010", 11795 => "10001000", 11796 => "01111101", 11802 => "10110000", 11806 => "11110101", 11807 => "00010011", 11809 => "00010111", 11813 => "11000111", 11814 => "11000101", 11815 => "10011101", 11816 => "10111101", 11818 => "10010110", 11820 => "11011001", 11821 => "00001100", 11822 => "01000011", 11823 => "01101000", 11826 => "01000011", 11829 => "01001000", 11833 => "10011111", 11834 => "10011111", 11835 => "11001111", 11836 => "01100000", 11837 => "00011010", 11838 => "10110110", 11839 => "00000100", 11841 => "10000011", 11842 => "01101001", 11844 => "10111011", 11845 => "11010000", 11846 => "01011101", 11847 => "11000111", 11848 => "00011010", 11852 => "00011000", 11853 => "01011111", 11855 => "01101100", 11856 => "11010010", 11857 => "10100100", 11858 => "10011111", 11859 => "01000110", 11860 => "10011101", 11862 => "11111000", 11864 => "11011111", 11865 => "01000100", 11866 => "01010111", 11868 => "11010111", 11869 => "10110010", 11870 => "00011001", 11871 => "10011000", 11872 => "00001100", 11875 => "10101110", 11879 => "01001101", 11880 => "01101100", 11881 => "00010100", 11883 => "00011101", 11888 => "10101110", 11889 => "01101100", 11890 => "00110000", 11892 => "10010111", 11894 => "10100111", 11896 => "01010011", 11898 => "01101001", 11899 => "01001101", 11900 => "00011110", 11901 => "10101111", 11903 => "00010001", 11904 => "01011111", 11905 => "01111010", 11907 => "00100000", 11908 => "01101000", 11911 => "10010011", 11913 => "10011110", 11914 => "10010011", 11915 => "00101010", 11917 => "00001011", 11918 => "00111101", 11919 => "11011011", 11920 => "01001010", 11921 => "11100001", 11922 => "01000111", 11929 => "11100000", 11934 => "11011010", 11935 => "10010010", 11936 => "00100010", 11938 => "10000001", 11941 => "10111010", 11942 => "00000110", 11946 => "01000011", 11948 => "10010100", 11950 => "10111001", 11953 => "10100111", 11954 => "00000011", 11955 => "00011101", 11956 => "11101111", 11959 => "00000100", 11960 => "00111110", 11961 => "11011111", 11962 => "01110100", 11963 => "01000101", 11965 => "00010000", 11967 => "01001011", 11968 => "01000011", 11973 => "10001011", 11974 => "10100010", 11976 => "10110000", 11977 => "11000000", 11978 => "11010011", 11979 => "11011111", 11985 => "11101010", 11986 => "11111001", 11988 => "11010000", 11992 => "01110100", 11995 => "00010101", 11996 => "00010000", 11999 => "00011110", 12003 => "10110010", 12004 => "00100010", 12005 => "00010110", 12008 => "11101111", 12009 => "10000000", 12013 => "11001111", 12015 => "11110110", 12016 => "10100100", 12020 => "10011110", 12022 => "01110000", 12023 => "11101000", 12029 => "01101011", 12030 => "10010010", 12032 => "11100100", 12034 => "11001011", 12036 => "01011011", 12040 => "10011110", 12042 => "01001000", 12043 => "00110010", 12044 => "01000010", 12046 => "01110111", 12048 => "10100010", 12052 => "00000100", 12062 => "10110110", 12064 => "10101101", 12065 => "10011100", 12066 => "11011100", 12068 => "10111110", 12069 => "00110111", 12073 => "01101100", 12075 => "11001011", 12077 => "01110101", 12078 => "11111000", 12079 => "01001110", 12083 => "10000010", 12085 => "00111000", 12086 => "01001101", 12090 => "10100101", 12092 => "10111000", 12095 => "01010101", 12096 => "11100010", 12098 => "10110001", 12099 => "01001111", 12101 => "10111011", 12103 => "11000110", 12104 => "01100101", 12108 => "00100000", 12118 => "00101011", 12123 => "00001110", 12126 => "01100100", 12127 => "10101101", 12128 => "11010101", 12133 => "01011100", 12136 => "11111001", 12139 => "01110110", 12140 => "11010110", 12141 => "11010101", 12142 => "10001011", 12144 => "10010110", 12147 => "11010100", 12151 => "01010110", 12152 => "11011111", 12153 => "00110100", 12154 => "00000100", 12156 => "01001010", 12159 => "10000010", 12161 => "01000111", 12163 => "00101010", 12164 => "01001010", 12166 => "01001001", 12171 => "01001101", 12172 => "00100101", 12174 => "11110100", 12175 => "11010010", 12176 => "00101000", 12180 => "11100011", 12186 => "01101000", 12187 => "10010001", 12189 => "01111101", 12190 => "00110111", 12194 => "01100101", 12196 => "01011111", 12202 => "00111011", 12205 => "10101011", 12206 => "00000001", 12207 => "11110111", 12209 => "01110101", 12211 => "00000010", 12212 => "11111001", 12214 => "10110000", 12215 => "10111101", 12219 => "10011000", 12224 => "11110011", 12229 => "01000000", 12230 => "10100111", 12231 => "00110011", 12234 => "01010110", 12235 => "00110000", 12237 => "11111000", 12239 => "00011000", 12241 => "00110101", 12244 => "01011000", 12245 => "00101111", 12246 => "00011110", 12247 => "11101111", 12250 => "11000100", 12251 => "10011001", 12256 => "00011010", 12257 => "10000000", 12261 => "01001010", 12262 => "01110101", 12265 => "00000111", 12266 => "00101101", 12267 => "11110101", 12268 => "00101100", 12272 => "00111100", 12278 => "01110111", 12279 => "11101100", 12280 => "11010100", 12281 => "00000101", 12282 => "10110111", 12283 => "01100110", 12284 => "11101000", 12287 => "10001101", 12288 => "11110101", 12289 => "11111110", 12290 => "01100111", 12292 => "10011101", 12293 => "11001110", 12296 => "01000001", 12298 => "11000111", 12300 => "11111110", 12302 => "01101001", 12304 => "11001111", 12308 => "10110111", 12310 => "11100000", 12311 => "10010111", 12312 => "11111011", 12314 => "00011010", 12315 => "11000011", 12316 => "10010011", 12321 => "01010000", 12323 => "00110011", 12324 => "00011001", 12325 => "11100001", 12327 => "00011001", 12328 => "01100001", 12329 => "01010011", 12332 => "10110000", 12333 => "11100100", 12335 => "01101100", 12336 => "10100001", 12337 => "11001111", 12338 => "01011111", 12339 => "11100100", 12340 => "11111110", 12341 => "11100011", 12344 => "01000111", 12345 => "00111000", 12346 => "11101101", 12349 => "01101101", 12352 => "00010100", 12355 => "10010011", 12356 => "01000101", 12357 => "11110011", 12362 => "10101100", 12370 => "00001111", 12371 => "01101011", 12373 => "10000110", 12375 => "00101001", 12376 => "10011010", 12379 => "01000001", 12381 => "00101100", 12385 => "01111111", 12394 => "01011001", 12397 => "11110100", 12399 => "10110100", 12400 => "01101111", 12402 => "10101011", 12405 => "01001000", 12407 => "10010111", 12408 => "01000110", 12409 => "10011001", 12411 => "01111010", 12413 => "01000000", 12415 => "11010111", 12416 => "11010100", 12417 => "01110110", 12418 => "10000001", 12421 => "10111000", 12422 => "01111111", 12424 => "11000000", 12426 => "11010110", 12430 => "01110001", 12431 => "11001000", 12434 => "01111011", 12437 => "10110110", 12442 => "01001010", 12445 => "00000111", 12447 => "01101110", 12453 => "01010011", 12454 => "10000000", 12455 => "11111011", 12456 => "10100100", 12457 => "10011111", 12458 => "11000010", 12459 => "01011101", 12460 => "10000100", 12462 => "00101001", 12463 => "10001010", 12464 => "11010111", 12466 => "11010010", 12467 => "10111011", 12468 => "11000001", 12469 => "10011101", 12470 => "10000101", 12471 => "11110101", 12472 => "00101001", 12473 => "10000100", 12478 => "01110110", 12480 => "11111110", 12482 => "01011100", 12486 => "10100011", 12490 => "11110001", 12493 => "01110010", 12496 => "01010110", 12498 => "01101011", 12499 => "00010111", 12500 => "11110111", 12501 => "11110110", 12503 => "10111100", 12504 => "11000010", 12505 => "01000000", 12507 => "01000010", 12508 => "11001001", 12509 => "00010110", 12511 => "10000111", 12514 => "00111001", 12521 => "11101011", 12522 => "10001000", 12524 => "10100011", 12528 => "00011100", 12529 => "00101100", 12530 => "01000110", 12531 => "10001000", 12533 => "10011001", 12536 => "01001000", 12537 => "00011110", 12539 => "01000101", 12540 => "11011111", 12541 => "10111101", 12543 => "00010111", 12544 => "00010010", 12547 => "00101100", 12550 => "01011001", 12551 => "11110000", 12554 => "01100000", 12555 => "10011001", 12559 => "00110101", 12560 => "01111110", 12563 => "00011111", 12565 => "00110100", 12572 => "10101000", 12573 => "00100010", 12574 => "11110011", 12578 => "01011010", 12579 => "11010011", 12580 => "11001110", 12582 => "10110110", 12583 => "11101010", 12584 => "10111010", 12585 => "10100011", 12587 => "10010011", 12588 => "10011011", 12594 => "10101011", 12596 => "10100101", 12601 => "01000101", 12603 => "10011010", 12604 => "00101010", 12605 => "00010111", 12606 => "11101110", 12607 => "10011000", 12609 => "00101000", 12610 => "10100001", 12615 => "11001010", 12620 => "00101110", 12623 => "10010101", 12624 => "10010111", 12625 => "10111100", 12626 => "10111001", 12627 => "10110101", 12628 => "11001100", 12630 => "10111110", 12634 => "11111111", 12636 => "11111111", 12637 => "11100000", 12638 => "11011110", 12640 => "01000100", 12645 => "01000011", 12651 => "00110000", 12653 => "00110111", 12654 => "01000101", 12657 => "11100111", 12660 => "01011100", 12661 => "11100111", 12662 => "11011100", 12672 => "01000001", 12673 => "01000111", 12674 => "10001010", 12675 => "10011101", 12678 => "11010010", 12680 => "10001101", 12681 => "01000111", 12682 => "10001001", 12685 => "10110101", 12687 => "10001110", 12688 => "01100111", 12690 => "01100100", 12693 => "01011010", 12695 => "00001011", 12697 => "01110001", 12701 => "10011011", 12703 => "00010110", 12705 => "00000101", 12706 => "10001000", 12708 => "10000000", 12710 => "00100001", 12711 => "00110100", 12713 => "00110011", 12714 => "11001000", 12719 => "00001001", 12721 => "10000000", 12722 => "11101101", 12726 => "00010100", 12727 => "11010000", 12734 => "11010011", 12735 => "00110100", 12737 => "11010010", 12739 => "11010111", 12741 => "10001001", 12743 => "01010001", 12748 => "01000010", 12751 => "10100001", 12753 => "00101110", 12755 => "01011111", 12756 => "01011110", 12758 => "00000100", 12760 => "01101011", 12762 => "10010000", 12763 => "11100110", 12766 => "00000100", 12769 => "11111110", 12771 => "00100001", 12774 => "00110000", 12775 => "00101111", 12781 => "01001110", 12783 => "01110011", 12784 => "10100111", 12785 => "00111111", 12788 => "10110100", 12789 => "00100111", 12794 => "11100011", 12795 => "11011011", 12796 => "01100011", 12797 => "10011000", 12798 => "00110100", 12800 => "00011010", 12806 => "00101111", 12808 => "01101100", 12810 => "01111111", 12811 => "00010001", 12820 => "01000101", 12822 => "11011000", 12824 => "10011110", 12832 => "10111111", 12835 => "10111110", 12837 => "00111100", 12841 => "01010001", 12842 => "10010010", 12849 => "01010001", 12851 => "00100110", 12856 => "00011011", 12864 => "10111110", 12866 => "01011000", 12880 => "11011000", 12881 => "10000000", 12884 => "11111110", 12885 => "10011101", 12886 => "01011010", 12887 => "10111010", 12888 => "00101111", 12889 => "11101011", 12890 => "10111000", 12891 => "00101101", 12893 => "11110101", 12897 => "00110001", 12902 => "10101100", 12906 => "01000000", 12907 => "10011100", 12910 => "11011000", 12911 => "00111000", 12912 => "11101111", 12913 => "01101010", 12915 => "00010000", 12916 => "11011001", 12919 => "11110101", 12920 => "10000111", 12922 => "11111101", 12923 => "00101110", 12927 => "11010011", 12928 => "11010110", 12932 => "01101001", 12933 => "00001100", 12935 => "10111010", 12936 => "10001110", 12937 => "10101000", 12946 => "01111100", 12947 => "01110000", 12951 => "10100101", 12953 => "11001111", 12954 => "10100001", 12956 => "01001001", 12959 => "10101011", 12960 => "11001011", 12966 => "00001011", 12967 => "01011010", 12970 => "00110001", 12972 => "10100101", 12973 => "10000111", 12979 => "01110010", 12981 => "10110101", 12984 => "11100100", 12985 => "01001000", 12986 => "00100101", 12987 => "10001110", 12988 => "01101111", 12990 => "10000010", 12991 => "11011101", 12992 => "10000101", 12993 => "00111011", 12995 => "01100100", 12998 => "00010011", 12999 => "10011100", 13000 => "11100011", 13003 => "00011110", 13005 => "01011000", 13008 => "00011101", 13014 => "00000111", 13015 => "11010101", 13017 => "10100111", 13021 => "11011001", 13022 => "11011010", 13023 => "10010101", 13025 => "11001010", 13028 => "01001010", 13029 => "01010100", 13030 => "10011101", 13031 => "10101100", 13032 => "00101010", 13034 => "00001111", 13037 => "00010010", 13045 => "10111101", 13046 => "11001011", 13047 => "01011000", 13049 => "00100000", 13052 => "00001001", 13053 => "11110100", 13054 => "11011100", 13055 => "11001101", 13058 => "10110111", 13062 => "10101111", 13065 => "10001111", 13066 => "11001000", 13067 => "11100011", 13070 => "11000110", 13071 => "01000111", 13074 => "01100001", 13079 => "11000100", 13082 => "00110100", 13084 => "11100010", 13086 => "00001111", 13092 => "11100110", 13096 => "11001001", 13100 => "10111000", 13101 => "11100011", 13102 => "01011101", 13103 => "10110101", 13104 => "11001100", 13105 => "10111000", 13106 => "01111011", 13109 => "01000101", 13110 => "01101011", 13116 => "01100100", 13118 => "11000111", 13119 => "11010110", 13120 => "11000000", 13125 => "00000110", 13127 => "11101000", 13128 => "11110100", 13135 => "11110010", 13136 => "11011111", 13138 => "11011010", 13140 => "01110101", 13141 => "01010100", 13142 => "11100111", 13143 => "01001111", 13144 => "01111001", 13145 => "10110000", 13146 => "01011001", 13148 => "11100000", 13150 => "11100100", 13152 => "00111111", 13154 => "11001110", 13157 => "00001100", 13162 => "00010110", 13166 => "10010011", 13169 => "00010101", 13171 => "11000100", 13172 => "00010100", 13173 => "10010111", 13175 => "11101011", 13177 => "10010001", 13179 => "01011110", 13181 => "11000111", 13183 => "00111101", 13186 => "01010010", 13189 => "00001101", 13191 => "10101111", 13192 => "10011110", 13200 => "11111101", 13203 => "00100001", 13204 => "00110100", 13207 => "10101110", 13208 => "01100011", 13211 => "01010101", 13212 => "11000111", 13213 => "10110110", 13215 => "01100011", 13218 => "01001011", 13220 => "11111011", 13224 => "11111110", 13226 => "00100100", 13228 => "11111100", 13230 => "00010011", 13231 => "10101100", 13233 => "10000111", 13234 => "10110100", 13235 => "10010110", 13236 => "01000000", 13237 => "10000101", 13243 => "10001001", 13244 => "01000000", 13247 => "00011110", 13249 => "11011101", 13251 => "10011111", 13252 => "11010010", 13253 => "01111111", 13255 => "01111001", 13256 => "00010100", 13258 => "11100100", 13261 => "10101111", 13262 => "01011000", 13264 => "10100000", 13267 => "01110001", 13268 => "11100101", 13269 => "11100111", 13270 => "00110010", 13271 => "11100110", 13272 => "10101010", 13277 => "10010011", 13279 => "10000101", 13280 => "01000001", 13281 => "00101011", 13282 => "01011110", 13283 => "10110011", 13284 => "11100010", 13286 => "01000100", 13287 => "01111101", 13289 => "01110000", 13294 => "10000100", 13296 => "10011110", 13298 => "10011010", 13299 => "11010000", 13300 => "00101001", 13302 => "11010110", 13304 => "00001010", 13306 => "00101110", 13308 => "00001110", 13311 => "10100010", 13314 => "00001001", 13315 => "00010011", 13316 => "01001110", 13317 => "00010100", 13321 => "10100011", 13322 => "10000000", 13325 => "01100100", 13326 => "10001010", 13330 => "11001011", 13332 => "01101001", 13333 => "10011000", 13335 => "11110100", 13340 => "11010101", 13342 => "00111111", 13344 => "01101000", 13346 => "01010100", 13348 => "10110110", 13349 => "11111111", 13351 => "10111100", 13354 => "11001111", 13355 => "10111111", 13357 => "10011100", 13360 => "00010100", 13361 => "10110001", 13362 => "01111011", 13368 => "11100001", 13372 => "11011110", 13375 => "11011010", 13377 => "00110111", 13378 => "10111101", 13379 => "11010110", 13384 => "10011000", 13386 => "01110100", 13387 => "00111001", 13388 => "00010111", 13392 => "00101101", 13395 => "01100011", 13397 => "01111000", 13400 => "10101010", 13401 => "01110110", 13402 => "01110010", 13404 => "00110000", 13407 => "10111110", 13409 => "01111001", 13410 => "00111111", 13411 => "01101010", 13412 => "01111010", 13413 => "01010110", 13414 => "11000111", 13416 => "11011010", 13417 => "01000100", 13418 => "01111011", 13425 => "10011011", 13426 => "11100110", 13427 => "11101000", 13428 => "01111101", 13429 => "01000001", 13430 => "10010000", 13434 => "00011011", 13436 => "00101000", 13444 => "00011100", 13445 => "01110000", 13449 => "01000101", 13450 => "00100000", 13456 => "11110111", 13457 => "00011101", 13458 => "01001000", 13459 => "01101111", 13461 => "10000001", 13465 => "10100110", 13470 => "11010000", 13471 => "10001010", 13472 => "01111010", 13473 => "00111010", 13478 => "01011100", 13480 => "00010110", 13482 => "10100000", 13484 => "01010000", 13487 => "10010101", 13488 => "11000000", 13490 => "01100011", 13491 => "01000010", 13493 => "01110100", 13496 => "00001100", 13499 => "00000010", 13500 => "00000001", 13501 => "01011001", 13502 => "00101111", 13503 => "11111110", 13504 => "00110010", 13506 => "10101111", 13507 => "10001100", 13509 => "01100011", 13511 => "00100000", 13513 => "11010101", 13514 => "01111010", 13515 => "01001011", 13516 => "01000011", 13517 => "01010010", 13520 => "11010101", 13521 => "10101101", 13522 => "11001110", 13527 => "01101101", 13533 => "11110111", 13534 => "11010000", 13535 => "00101100", 13536 => "01000001", 13537 => "01011001", 13538 => "00010011", 13539 => "00000010", 13541 => "11011010", 13544 => "10110100", 13546 => "10010101", 13548 => "11101110", 13550 => "00010110", 13553 => "11001100", 13554 => "10101111", 13555 => "00010110", 13557 => "11001010", 13558 => "01011000", 13559 => "10101000", 13560 => "00010110", 13564 => "01111000", 13565 => "10111011", 13569 => "11111101", 13570 => "11000101", 13571 => "10010000", 13572 => "10110100", 13574 => "11111011", 13575 => "11000100", 13578 => "11100101", 13579 => "01101101", 13580 => "10100111", 13581 => "00000010", 13582 => "11111000", 13583 => "01100111", 13586 => "01101011", 13590 => "10111011", 13592 => "10011001", 13594 => "11001011", 13595 => "10100110", 13597 => "00010111", 13598 => "11100111", 13601 => "11010110", 13610 => "10100010", 13611 => "00011011", 13613 => "11010111", 13614 => "11001111", 13615 => "00010100", 13616 => "11101101", 13618 => "11111101", 13623 => "11100001", 13626 => "01000011", 13627 => "00000101", 13629 => "11010011", 13630 => "11111110", 13631 => "01100001", 13634 => "01011010", 13638 => "11101010", 13639 => "11110010", 13640 => "01100001", 13641 => "11011001", 13644 => "00110001", 13646 => "01011100", 13648 => "10001110", 13649 => "01010101", 13651 => "10010000", 13652 => "11101000", 13653 => "10100111", 13656 => "01101110", 13660 => "11010010", 13663 => "01011100", 13664 => "01100000", 13668 => "10111000", 13670 => "01101001", 13675 => "11001010", 13677 => "00001010", 13679 => "01100010", 13680 => "01100010", 13681 => "00000100", 13682 => "00010011", 13685 => "10011100", 13688 => "00011011", 13689 => "10101010", 13694 => "10110100", 13696 => "11111111", 13697 => "10111110", 13701 => "01110011", 13702 => "10000100", 13705 => "11100110", 13706 => "00100001", 13707 => "11000001", 13711 => "10010101", 13715 => "10001111", 13716 => "10111100", 13717 => "00010101", 13718 => "10100100", 13722 => "01001111", 13725 => "01010110", 13727 => "11010000", 13729 => "00100101", 13730 => "10110011", 13731 => "01100001", 13733 => "10000111", 13736 => "11110101", 13739 => "00100010", 13740 => "10100101", 13741 => "10111101", 13742 => "01000110", 13746 => "01101011", 13747 => "01001001", 13748 => "00011011", 13749 => "10111001", 13750 => "10000011", 13751 => "01001100", 13752 => "01000110", 13753 => "01111001", 13754 => "00001001", 13755 => "01110010", 13756 => "01101110", 13761 => "01010000", 13763 => "11010110", 13765 => "01011110", 13767 => "11001111", 13768 => "11111001", 13771 => "10001110", 13772 => "11011101", 13774 => "01111010", 13777 => "10000000", 13778 => "00101010", 13782 => "01101110", 13790 => "01100011", 13792 => "11100010", 13794 => "10110111", 13798 => "11101011", 13801 => "00001011", 13802 => "10111001", 13805 => "10111100", 13806 => "01111010", 13808 => "11001101", 13809 => "00001101", 13811 => "11110111", 13813 => "01001001", 13815 => "10001100", 13818 => "11010001", 13819 => "01101011", 13820 => "11101001", 13821 => "11000001", 13822 => "10001110", 13823 => "11101011", 13824 => "11001011", 13825 => "01111000", 13827 => "11011110", 13831 => "10001110", 13832 => "01110110", 13833 => "00001100", 13834 => "10011001", 13836 => "00110010", 13837 => "11011010", 13838 => "00001011", 13840 => "00110100", 13845 => "11010110", 13847 => "00100001", 13848 => "01010101", 13849 => "10001011", 13851 => "01111000", 13852 => "01100110", 13860 => "00110110", 13861 => "11001001", 13864 => "10111010", 13866 => "00101110", 13868 => "11100110", 13870 => "10010101", 13873 => "11100100", 13877 => "01000010", 13878 => "11001110", 13880 => "10110101", 13881 => "11010111", 13882 => "11000000", 13883 => "11100000", 13886 => "11000101", 13890 => "01110100", 13892 => "10000001", 13893 => "01110100", 13898 => "01101011", 13903 => "01001011", 13905 => "11011110", 13908 => "00001110", 13909 => "01100011", 13912 => "00011111", 13920 => "10010101", 13923 => "11111000", 13925 => "10100010", 13926 => "01001010", 13930 => "11100111", 13931 => "10000110", 13935 => "11110000", 13938 => "00101001", 13939 => "11110100", 13943 => "00111001", 13944 => "10011011", 13946 => "00100110", 13947 => "11101101", 13948 => "00001100", 13950 => "10000100", 13951 => "10000110", 13952 => "01100011", 13953 => "10011001", 13954 => "11000011", 13956 => "00111010", 13959 => "01000001", 13964 => "10110001", 13970 => "00110111", 13971 => "11000010", 13972 => "00111000", 13973 => "01001110", 13974 => "10001010", 13976 => "01111100", 13978 => "00101101", 13980 => "00001010", 13981 => "00110011", 13982 => "00001110", 13983 => "10001010", 13985 => "01000010", 13990 => "10101100", 13991 => "00100100", 13993 => "00011010", 13994 => "00000110", 13995 => "01011100", 13996 => "01111011", 13997 => "01011000", 13999 => "00101110", 14001 => "11010001", 14002 => "00000111", 14004 => "11111001", 14007 => "00011111", 14011 => "00101110", 14012 => "10110010", 14017 => "00011101", 14018 => "11110101", 14020 => "00110010", 14023 => "11111010", 14025 => "01101000", 14030 => "10000001", 14032 => "01000101", 14036 => "00100000", 14037 => "00100100", 14039 => "11100011", 14040 => "01111001", 14043 => "01101100", 14045 => "01101100", 14046 => "01000000", 14049 => "11010011", 14050 => "00000100", 14052 => "00110001", 14053 => "11011011", 14059 => "10101000", 14060 => "01000100", 14064 => "10110000", 14066 => "01001110", 14067 => "11011011", 14070 => "11010100", 14077 => "10001101", 14080 => "11100001", 14081 => "01000010", 14082 => "11010000", 14085 => "11100011", 14086 => "11001000", 14090 => "10010000", 14091 => "10010010", 14095 => "10001100", 14096 => "01111100", 14097 => "00010110", 14098 => "01101011", 14099 => "11010110", 14100 => "00100110", 14101 => "11101000", 14107 => "00110000", 14109 => "00110101", 14110 => "11010101", 14112 => "11001111", 14116 => "10110010", 14117 => "00000110", 14120 => "10010110", 14121 => "10101011", 14122 => "10101011", 14124 => "11110101", 14126 => "00011011", 14127 => "11110110", 14129 => "10100001", 14130 => "11101101", 14132 => "00101100", 14133 => "00001100", 14134 => "01011000", 14135 => "00111010", 14136 => "11110011", 14137 => "10011011", 14139 => "01101000", 14142 => "00101101", 14143 => "10100001", 14146 => "11101110", 14152 => "00000011", 14155 => "10000110", 14156 => "10001110", 14157 => "01111011", 14158 => "10000011", 14159 => "10010010", 14160 => "01111001", 14162 => "11010100", 14164 => "11101111", 14165 => "10001101", 14166 => "11111111", 14170 => "11000011", 14171 => "00110110", 14172 => "10001100", 14174 => "00110111", 14175 => "00011110", 14177 => "01100111", 14180 => "00010010", 14188 => "00100000", 14189 => "11110101", 14193 => "10011000", 14196 => "10100111", 14197 => "00011000", 14199 => "01000001", 14200 => "11000001", 14202 => "01011000", 14203 => "11001011", 14204 => "00011110", 14208 => "01100101", 14210 => "00000011", 14214 => "11001001", 14215 => "00001010", 14221 => "00100110", 14222 => "01011011", 14225 => "01010100", 14226 => "11110101", 14228 => "11111110", 14229 => "01001110", 14231 => "10011110", 14232 => "01010011", 14233 => "11011001", 14234 => "10001001", 14235 => "11111011", 14236 => "01101110", 14237 => "11111011", 14242 => "01110001", 14243 => "10011011", 14245 => "01110010", 14248 => "00001101", 14249 => "01000011", 14251 => "10101101", 14255 => "10101110", 14257 => "01100100", 14259 => "10010101", 14260 => "11110111", 14262 => "01100000", 14264 => "00011100", 14266 => "11001010", 14269 => "11010110", 14271 => "10110100", 14272 => "01010011", 14274 => "01111100", 14275 => "11010101", 14277 => "11101010", 14278 => "11100001", 14283 => "00111000", 14285 => "00111101", 14287 => "11111001", 14288 => "01000101", 14291 => "01000101", 14292 => "00111011", 14293 => "10110010", 14295 => "10000111", 14298 => "10111111", 14302 => "10100011", 14303 => "00101000", 14305 => "01100011", 14306 => "11000111", 14307 => "00110000", 14308 => "00101100", 14309 => "10111100", 14310 => "11010000", 14311 => "01011011", 14312 => "11001101", 14313 => "10110001", 14315 => "00001011", 14319 => "01110010", 14321 => "10110010", 14322 => "10110000", 14325 => "00000001", 14326 => "00001110", 14327 => "11010100", 14328 => "10011010", 14329 => "11011000", 14331 => "10011000", 14332 => "01000101", 14333 => "10011001", 14334 => "11101111", 14336 => "11101011", 14337 => "01000101", 14339 => "11011110", 14340 => "01110100", 14341 => "11111100", 14342 => "10010100", 14343 => "11010100", 14345 => "10001010", 14353 => "11000100", 14354 => "10010110", 14358 => "10100101", 14359 => "11000010", 14360 => "01010100", 14362 => "00110110", 14363 => "10101001", 14364 => "10100000", 14367 => "10101111", 14369 => "00001111", 14372 => "10010001", 14374 => "10000111", 14376 => "11000011", 14378 => "11001011", 14380 => "11010101", 14388 => "11000001", 14389 => "01010110", 14390 => "00010101", 14392 => "11101111", 14393 => "00101110", 14394 => "11101100", 14395 => "11000110", 14397 => "11001111", 14398 => "10010000", 14399 => "10100100", 14402 => "10001010", 14403 => "10001100", 14404 => "11000010", 14405 => "11001001", 14407 => "11110000", 14409 => "01110000", 14410 => "10110100", 14411 => "00011101", 14413 => "11001000", 14414 => "00011101", 14417 => "11110101", 14418 => "10110101", 14419 => "10100110", 14423 => "11001100", 14424 => "01010001", 14425 => "01101110", 14427 => "01010000", 14431 => "11101000", 14432 => "10111111", 14433 => "11101010", 14435 => "11101100", 14438 => "10101101", 14440 => "11110000", 14441 => "00000111", 14443 => "11101001", 14446 => "10001100", 14448 => "00011010", 14453 => "11010011", 14455 => "11110011", 14456 => "11000011", 14458 => "11111011", 14459 => "00010000", 14462 => "10010001", 14464 => "10101101", 14466 => "00010101", 14470 => "10110001", 14471 => "11110000", 14473 => "00100010", 14474 => "11010010", 14475 => "11111000", 14477 => "10001100", 14483 => "11101010", 14485 => "00000011", 14486 => "00100110", 14489 => "00100111", 14490 => "11000101", 14495 => "01001011", 14497 => "00101011", 14502 => "01001110", 14503 => "11000110", 14507 => "10110110", 14509 => "10111110", 14518 => "00001111", 14520 => "11100000", 14521 => "01001110", 14523 => "10110111", 14524 => "01010111", 14525 => "00010000", 14530 => "01011001", 14533 => "11011111", 14534 => "11010101", 14536 => "10010101", 14538 => "01011010", 14539 => "10001001", 14541 => "01101001", 14542 => "00001110", 14543 => "10100001", 14546 => "00011111", 14549 => "10010010", 14552 => "10110011", 14553 => "11101011", 14555 => "00011000", 14556 => "10110010", 14558 => "01111000", 14560 => "01100010", 14561 => "00000101", 14562 => "11110111", 14563 => "11000100", 14564 => "11001000", 14569 => "11000001", 14570 => "00101000", 14572 => "00011110", 14575 => "10110110", 14578 => "10001111", 14581 => "10001010", 14583 => "00011111", 14584 => "10111111", 14585 => "11100011", 14586 => "11100101", 14587 => "11101010", 14588 => "00110101", 14591 => "00010010", 14593 => "10010010", 14595 => "10011001", 14597 => "01011011", 14602 => "01111111", 14604 => "10101011", 14608 => "10100101", 14609 => "00001111", 14610 => "01001000", 14612 => "10110011", 14613 => "00000001", 14616 => "11000000", 14618 => "11110111", 14619 => "11001100", 14621 => "10111101", 14624 => "10101000", 14625 => "00101110", 14627 => "10111001", 14628 => "11110001", 14629 => "11010111", 14630 => "11010011", 14631 => "10101010", 14636 => "00001110", 14637 => "10011101", 14638 => "00001111", 14639 => "10100111", 14641 => "10101100", 14642 => "01111011", 14643 => "11100110", 14645 => "11000110", 14647 => "10011011", 14648 => "01001010", 14649 => "11101101", 14650 => "11110001", 14651 => "00011011", 14652 => "01010100", 14653 => "10011101", 14654 => "00001010", 14656 => "10011011", 14657 => "01111110", 14658 => "00100101", 14659 => "01011010", 14660 => "00101111", 14663 => "01101011", 14670 => "11111101", 14671 => "11111110", 14675 => "10010000", 14676 => "11111101", 14678 => "10100001", 14683 => "01111111", 14684 => "00110011", 14685 => "11100110", 14694 => "00101001", 14695 => "01010001", 14697 => "11011011", 14698 => "01010111", 14699 => "10000010", 14700 => "00100110", 14701 => "01010001", 14707 => "01000011", 14708 => "10011010", 14711 => "00011100", 14714 => "00010110", 14715 => "01010111", 14716 => "11000011", 14717 => "10001010", 14722 => "11000001", 14724 => "11110000", 14726 => "10000001", 14731 => "11011011", 14734 => "01100100", 14735 => "01001111", 14737 => "00000010", 14738 => "10111001", 14739 => "01100110", 14746 => "00011100", 14747 => "01111011", 14748 => "00110010", 14752 => "11011111", 14757 => "10111001", 14758 => "10111101", 14761 => "00101110", 14770 => "01100110", 14771 => "01010001", 14773 => "11011100", 14774 => "11101010", 14775 => "00110010", 14781 => "00001110", 14786 => "10110010", 14787 => "01111011", 14789 => "11100101", 14791 => "11111001", 14792 => "10101000", 14793 => "10111111", 14794 => "00001111", 14795 => "00011011", 14796 => "11010110", 14800 => "11000111", 14802 => "11000111", 14803 => "11001001", 14809 => "10001111", 14813 => "01000000", 14815 => "00010010", 14816 => "01010100", 14817 => "00110011", 14818 => "01001010", 14819 => "10100100", 14824 => "01011100", 14825 => "11111000", 14826 => "01000101", 14829 => "11000001", 14833 => "11110011", 14835 => "01000111", 14837 => "11010001", 14839 => "00000001", 14842 => "11000101", 14843 => "01100110", 14845 => "11110011", 14848 => "10010011", 14849 => "00100000", 14850 => "10001001", 14851 => "01001011", 14855 => "00000111", 14858 => "10001100", 14860 => "01010001", 14864 => "11100000", 14866 => "11010000", 14867 => "01100110", 14868 => "01101010", 14870 => "01000111", 14872 => "11000101", 14873 => "01100110", 14874 => "01100000", 14876 => "11010001", 14877 => "00111111", 14879 => "10001101", 14880 => "01111101", 14881 => "11011111", 14883 => "01110111", 14884 => "00101100", 14886 => "00001111", 14887 => "01111001", 14888 => "00010000", 14889 => "01001111", 14890 => "11010100", 14892 => "01010110", 14893 => "11000000", 14896 => "00010100", 14897 => "01111111", 14899 => "00100101", 14900 => "10011001", 14906 => "00001111", 14907 => "10001001", 14909 => "10001100", 14912 => "00100111", 14914 => "00111111", 14916 => "01011111", 14920 => "01001001", 14922 => "11100001", 14923 => "00011100", 14924 => "01111001", 14927 => "01110101", 14928 => "00111001", 14929 => "10011011", 14930 => "10000100", 14934 => "10001001", 14935 => "11101110", 14937 => "10000001", 14939 => "01011011", 14942 => "00101101", 14943 => "01001101", 14944 => "10000011", 14950 => "00110000", 14952 => "11001000", 14953 => "01101001", 14958 => "10110010", 14959 => "01100011", 14960 => "00111101", 14961 => "11100001", 14962 => "11100001", 14963 => "11100100", 14967 => "01101110", 14968 => "11001000", 14970 => "11011011", 14971 => "01011000", 14974 => "11010110", 14975 => "10100011", 14976 => "01111001", 14978 => "00000101", 14981 => "10100101", 14983 => "10001011", 14986 => "00000101", 14987 => "01111000", 14990 => "11100010", 14993 => "10111110", 14994 => "10111111", 14995 => "10000101", 14997 => "11001011", 14999 => "11100011", 15002 => "11011000", 15006 => "10101101", 15007 => "01100011", 15009 => "11001001", 15010 => "00101101", 15011 => "00000001", 15012 => "11110111", 15015 => "11110010", 15016 => "00110100", 15022 => "11011100", 15024 => "00111011", 15027 => "00001011", 15029 => "01010101", 15030 => "10001001", 15031 => "11001000", 15033 => "10101011", 15034 => "01000100", 15035 => "00010011", 15037 => "01011110", 15041 => "01101001", 15043 => "10100001", 15045 => "01101010", 15046 => "01100000", 15048 => "01001100", 15051 => "11011010", 15052 => "11100001", 15056 => "10001010", 15057 => "01101010", 15058 => "01000001", 15059 => "00010010", 15060 => "10010011", 15067 => "01100001", 15068 => "00101000", 15069 => "10010000", 15071 => "00011100", 15073 => "00010011", 15076 => "10101000", 15077 => "00101000", 15079 => "00101111", 15080 => "00001101", 15082 => "00011111", 15083 => "11101011", 15086 => "00000001", 15091 => "01011111", 15094 => "11011110", 15095 => "00000001", 15096 => "00010100", 15098 => "00110111", 15100 => "10110001", 15101 => "11001111", 15102 => "01101010", 15103 => "11110011", 15106 => "11101101", 15107 => "11110000", 15109 => "11011000", 15110 => "00110100", 15111 => "10000100", 15112 => "11011001", 15119 => "10001110", 15123 => "10110111", 15126 => "10110100", 15129 => "01101010", 15130 => "00101101", 15132 => "00110000", 15136 => "00110001", 15137 => "11101001", 15139 => "10101011", 15140 => "00100111", 15142 => "00001011", 15144 => "11011010", 15146 => "11001101", 15149 => "11101000", 15150 => "00110000", 15152 => "11100010", 15153 => "10000101", 15155 => "10001100", 15156 => "00110001", 15157 => "11110100", 15158 => "01101000", 15159 => "00000010", 15161 => "01001110", 15164 => "01101000", 15167 => "01111110", 15168 => "01111110", 15170 => "01100010", 15171 => "10100101", 15176 => "10101010", 15178 => "10010011", 15179 => "10001101", 15183 => "11110011", 15186 => "00100100", 15189 => "00011000", 15191 => "00101100", 15192 => "10101111", 15193 => "01100100", 15194 => "01010000", 15196 => "11001000", 15199 => "11110101", 15200 => "11001000", 15201 => "00101010", 15202 => "00110100", 15203 => "10110011", 15205 => "10111010", 15206 => "10000101", 15209 => "01000100", 15211 => "01110110", 15213 => "01110011", 15214 => "00101100", 15217 => "10010111", 15218 => "10100100", 15223 => "10101000", 15224 => "00111111", 15226 => "11000010", 15230 => "01101001", 15231 => "01101101", 15233 => "01011011", 15235 => "01101110", 15239 => "00111100", 15242 => "11101100", 15243 => "10100000", 15246 => "11010001", 15247 => "10101110", 15248 => "00011001", 15249 => "11110000", 15250 => "11001000", 15251 => "00001000", 15254 => "10001000", 15255 => "10101111", 15259 => "00101010", 15260 => "11001100", 15263 => "00100111", 15265 => "11101110", 15267 => "00111010", 15268 => "00001100", 15270 => "10100101", 15272 => "01101100", 15274 => "01111110", 15275 => "10001110", 15276 => "11111011", 15277 => "10001001", 15278 => "10101100", 15281 => "11111110", 15284 => "11001100", 15285 => "00011011", 15286 => "10110111", 15287 => "01001010", 15288 => "00001101", 15290 => "10000011", 15303 => "01001001", 15304 => "10001011", 15305 => "00110011", 15306 => "10011001", 15309 => "01011110", 15311 => "11110010", 15312 => "11100101", 15317 => "00010011", 15318 => "10111100", 15319 => "11100110", 15320 => "11011001", 15321 => "10111101", 15323 => "00110111", 15331 => "11110000", 15333 => "10011011", 15336 => "10101111", 15337 => "10100010", 15340 => "00010010", 15341 => "01110111", 15343 => "10100001", 15346 => "11111000", 15348 => "00001110", 15349 => "00011000", 15351 => "01101100", 15355 => "01010101", 15359 => "11001011", 15362 => "00000110", 15363 => "01010010", 15364 => "11010110", 15370 => "11100110", 15371 => "10000001", 15374 => "01001000", 15376 => "11000000", 15377 => "11100011", 15379 => "11011110", 15380 => "00011011", 15382 => "10101101", 15384 => "00110010", 15391 => "10111101", 15392 => "01000111", 15393 => "11100000", 15394 => "00010100", 15395 => "11110001", 15396 => "01100111", 15397 => "10110110", 15399 => "01101001", 15403 => "11011110", 15408 => "01001011", 15409 => "10100111", 15410 => "10010100", 15412 => "00010101", 15413 => "01000100", 15415 => "01000110", 15417 => "11010101", 15418 => "01100111", 15419 => "01111000", 15424 => "00110010", 15427 => "10110110", 15429 => "11101100", 15430 => "11111001", 15432 => "10101100", 15433 => "11010011", 15435 => "10001111", 15439 => "00000010", 15440 => "00010001", 15443 => "01000010", 15450 => "10111010", 15451 => "11011101", 15455 => "00011111", 15457 => "10110101", 15460 => "11111110", 15462 => "10110001", 15463 => "10010111", 15464 => "11101100", 15466 => "11100101", 15467 => "00010100", 15469 => "11101011", 15470 => "11010011", 15471 => "11001111", 15472 => "10100000", 15477 => "10000110", 15478 => "00100110", 15480 => "11101011", 15481 => "01001111", 15483 => "10111110", 15484 => "00101101", 15488 => "10011001", 15489 => "11111001", 15494 => "10000011", 15495 => "11000111", 15498 => "00111100", 15499 => "00100000", 15501 => "11100100", 15502 => "10110101", 15503 => "00001101", 15504 => "11000001", 15507 => "00110111", 15513 => "01110111", 15516 => "01011111", 15518 => "10001110", 15519 => "00110010", 15520 => "10010111", 15522 => "10110010", 15523 => "10011001", 15525 => "11001000", 15533 => "11111110", 15534 => "11111001", 15536 => "01000100", 15537 => "01111100", 15538 => "10011110", 15541 => "01100011", 15542 => "11111000", 15545 => "00111110", 15547 => "00010000", 15552 => "11100101", 15554 => "10111101", 15555 => "11000111", 15556 => "11100011", 15557 => "11000010", 15560 => "01010111", 15562 => "10010011", 15567 => "11101111", 15568 => "10100000", 15570 => "10001100", 15571 => "10110101", 15574 => "00001101", 15577 => "01000110", 15579 => "10110110", 15580 => "11100110", 15583 => "00100111", 15584 => "11011111", 15586 => "11001011", 15587 => "00001100", 15588 => "11101001", 15589 => "10101011", 15591 => "10101100", 15592 => "10011001", 15594 => "10001101", 15595 => "11011010", 15596 => "10110111", 15597 => "11000001", 15599 => "01000110", 15600 => "11111001", 15601 => "00110001", 15602 => "01010101", 15603 => "10101010", 15606 => "10010111", 15607 => "10010001", 15611 => "00010001", 15612 => "10010100", 15613 => "10100001", 15614 => "11100010", 15617 => "10111100", 15619 => "11110110", 15620 => "11101110", 15622 => "01111011", 15624 => "11001011", 15625 => "10001100", 15627 => "10010000", 15628 => "01100110", 15629 => "00000101", 15630 => "10101010", 15631 => "00110011", 15637 => "10001001", 15639 => "11100110", 15640 => "01001001", 15642 => "01111010", 15645 => "11100010", 15646 => "00110110", 15650 => "11110100", 15651 => "01100010", 15652 => "10110011", 15653 => "11100001", 15654 => "00101010", 15658 => "01011011", 15661 => "00010011", 15664 => "10000000", 15666 => "00001101", 15667 => "11110000", 15671 => "00011001", 15673 => "01010010", 15674 => "10110111", 15677 => "00010010", 15679 => "00100111", 15680 => "00011100", 15682 => "01100000", 15684 => "00000010", 15686 => "11000100", 15687 => "11101011", 15692 => "11011111", 15693 => "11101101", 15696 => "00100110", 15697 => "11100110", 15700 => "11111000", 15703 => "11001100", 15706 => "11000100", 15707 => "01111011", 15710 => "00100111", 15713 => "10100110", 15714 => "01101000", 15715 => "01100101", 15716 => "10110100", 15717 => "01100100", 15718 => "01010101", 15721 => "10101101", 15728 => "00100000", 15730 => "11101100", 15731 => "11001110", 15733 => "01101101", 15736 => "11010100", 15741 => "00001110", 15743 => "01110100", 15744 => "10110011", 15745 => "11100110", 15749 => "10101111", 15750 => "11110101", 15753 => "00101010", 15756 => "00111111", 15757 => "00101110", 15758 => "00111111", 15760 => "00111111", 15762 => "10111100", 15766 => "00011101", 15770 => "01110010", 15771 => "10010011", 15772 => "11101110", 15773 => "11110010", 15774 => "00111101", 15777 => "01001011", 15778 => "10011111", 15780 => "01101111", 15787 => "00011110", 15788 => "11101010", 15789 => "01001100", 15791 => "10110001", 15793 => "00011110", 15796 => "10010000", 15797 => "01100111", 15799 => "10010011", 15801 => "10001100", 15802 => "00111001", 15804 => "11110101", 15818 => "01100100", 15820 => "01111000", 15821 => "01111100", 15822 => "10110000", 15825 => "11101100", 15827 => "10110101", 15829 => "10101110", 15831 => "11111101", 15832 => "01011011", 15833 => "11011011", 15837 => "01010100", 15838 => "10100110", 15842 => "10011001", 15844 => "11001110", 15845 => "01000000", 15847 => "11100101", 15849 => "10011111", 15850 => "00001010", 15851 => "00110111", 15857 => "01100111", 15862 => "11011000", 15863 => "00010001", 15866 => "00000111", 15868 => "10111111", 15872 => "11000000", 15874 => "01100111", 15876 => "11111100", 15878 => "11100011", 15880 => "11101000", 15881 => "01100110", 15883 => "00101101", 15886 => "10100110", 15888 => "00010100", 15889 => "00000100", 15891 => "01101001", 15893 => "10001010", 15896 => "10001001", 15897 => "11111100", 15898 => "11111100", 15900 => "11100101", 15903 => "00010111", 15906 => "11000011", 15912 => "11111110", 15914 => "11110000", 15918 => "01101000", 15919 => "00100111", 15927 => "10100101", 15932 => "01000111", 15933 => "00001100", 15934 => "11010011", 15935 => "10010010", 15937 => "01011110", 15939 => "00001000", 15940 => "10010000", 15941 => "11101110", 15944 => "10100010", 15950 => "00001011", 15952 => "11100101", 15953 => "00010100", 15955 => "11111011", 15958 => "01001011", 15959 => "10010011", 15960 => "00000110", 15961 => "11100011", 15965 => "01001110", 15972 => "10000010", 15974 => "10000000", 15977 => "11111101", 15981 => "00010000", 15982 => "10101101", 15986 => "00001000", 15989 => "11011011", 15991 => "00110110", 15993 => "01001011", 15996 => "10011010", 15997 => "01111000", 15999 => "00101101", 16000 => "10100110", 16004 => "11110111", 16009 => "00100001", 16010 => "01000101", 16011 => "11010011", 16014 => "11111101", 16017 => "10101011", 16018 => "11111110", 16019 => "00100110", 16020 => "00100011", 16021 => "11101110", 16022 => "00110001", 16024 => "00100001", 16026 => "00111111", 16028 => "10100110", 16030 => "01101011", 16034 => "11101010", 16036 => "01010000", 16041 => "00001110", 16044 => "01100011", 16045 => "00010100", 16046 => "10010111", 16047 => "01100000", 16048 => "00111100", 16054 => "11001111", 16055 => "11111111", 16056 => "11100010", 16057 => "11001001", 16058 => "11000101", 16059 => "01010001", 16061 => "11111101", 16063 => "11101010", 16064 => "11000010", 16065 => "01101101", 16066 => "11110101", 16070 => "00110101", 16071 => "11011011", 16073 => "11110000", 16074 => "11000100", 16076 => "00011011", 16080 => "00101000", 16081 => "00111001", 16085 => "00101010", 16087 => "10001111", 16089 => "01110101", 16093 => "10101111", 16094 => "10010000", 16095 => "01001100", 16099 => "00010100", 16105 => "00101001", 16106 => "01001110", 16110 => "10111100", 16112 => "10111001", 16113 => "00111111", 16114 => "01000001", 16117 => "00110011", 16120 => "10011100", 16121 => "10011111", 16122 => "01100011", 16124 => "00000010", 16127 => "00010001", 16128 => "00011111", 16129 => "10011010", 16131 => "10001000", 16132 => "01101011", 16133 => "10010101", 16135 => "00110011", 16138 => "11010111", 16139 => "01011011", 16141 => "11010010", 16142 => "00011111", 16143 => "11000011", 16144 => "11000000", 16147 => "10101011", 16149 => "10110000", 16150 => "00100010", 16151 => "10001000", 16155 => "10000000", 16157 => "01011001", 16158 => "10100111", 16162 => "01110101", 16165 => "01110100", 16167 => "01110100", 16168 => "01101010", 16173 => "11110001", 16178 => "00000010", 16181 => "10111001", 16182 => "11110101", 16184 => "01101000", 16186 => "10111110", 16188 => "10001110", 16189 => "11000001", 16193 => "00100101", 16195 => "00101010", 16196 => "00001000", 16197 => "10110101", 16198 => "00110010", 16201 => "01111100", 16202 => "01001100", 16204 => "10101011", 16207 => "01011101", 16210 => "00010110", 16211 => "11101110", 16213 => "01001111", 16215 => "10111111", 16217 => "10110111", 16220 => "11111011", 16221 => "10010011", 16223 => "00000001", 16225 => "10101010", 16227 => "11100000", 16229 => "10011011", 16230 => "00101101", 16231 => "11110110", 16233 => "10000000", 16234 => "10000010", 16235 => "10110111", 16237 => "10101011", 16239 => "11011000", 16242 => "01011111", 16244 => "11110100", 16247 => "11000110", 16248 => "10000011", 16249 => "01111101", 16250 => "01111010", 16251 => "01110001", 16252 => "11111010", 16255 => "10011001", 16256 => "00111111", 16260 => "00010000", 16263 => "11110100", 16264 => "10111110", 16265 => "10100011", 16269 => "01011111", 16273 => "10010000", 16274 => "11010000", 16276 => "11001110", 16277 => "01100001", 16279 => "11010001", 16280 => "11000100", 16282 => "00110110", 16286 => "00100011", 16287 => "01000100", 16290 => "11100000", 16292 => "11111101", 16293 => "01000110", 16294 => "00010000", 16296 => "01110000", 16298 => "00001011", 16300 => "00111011", 16301 => "01000000", 16303 => "00001011", 16308 => "01011100", 16309 => "00000001", 16310 => "01001110", 16311 => "01100000", 16312 => "10101010", 16315 => "00100111", 16317 => "10010000", 16320 => "01011110", 16322 => "10111101", 16326 => "00010100", 16327 => "00100101", 16330 => "10101011", 16331 => "11010101", 16336 => "00100011", 16338 => "00010110", 16339 => "01110110", 16343 => "10001101", 16346 => "01000011", 16353 => "00100101", 16356 => "11100011", 16358 => "01101010", 16362 => "10001110", 16363 => "11000001", 16366 => "00100010", 16367 => "01011011", 16369 => "11101100", 16376 => "10111011", 16377 => "01001011", 16379 => "10111010", 16380 => "01110000", 16382 => "00011110", 16385 => "11000100", 16388 => "11001110", 16390 => "00011101", 16394 => "10111011", 16395 => "11011010", 16398 => "01001011", 16399 => "11100110", 16401 => "00011101", 16402 => "01001111", 16403 => "01111001", 16410 => "00000101", 16412 => "10011110", 16413 => "01010011", 16416 => "00101100", 16420 => "00111110", 16430 => "01001101", 16431 => "01111000", 16435 => "10101101", 16437 => "10010001", 16439 => "00101111", 16442 => "00010000", 16443 => "01111101", 16445 => "10100000", 16448 => "01000111", 16449 => "10111010", 16450 => "11001101", 16456 => "10101010", 16457 => "01000010", 16458 => "11011010", 16459 => "01100101", 16461 => "11000000", 16462 => "11100010", 16464 => "01001011", 16465 => "10001000", 16467 => "01111110", 16468 => "01011001", 16469 => "01101101", 16471 => "00110110", 16477 => "01011001", 16479 => "00100010", 16480 => "01000100", 16481 => "01010111", 16483 => "01101101", 16484 => "10000110", 16485 => "00001111", 16486 => "11000111", 16489 => "01100001", 16490 => "01100110", 16491 => "01110110", 16493 => "00001101", 16495 => "01001100", 16496 => "10100100", 16498 => "00010010", 16501 => "10110011", 16502 => "01011010", 16503 => "11101000", 16505 => "10000001", 16506 => "01111110", 16507 => "11101111", 16508 => "01000001", 16509 => "01000100", 16513 => "01101000", 16514 => "00010001", 16516 => "10111100", 16517 => "10110001", 16519 => "10111101", 16522 => "00111011", 16524 => "10100001", 16525 => "00100111", 16526 => "10111011", 16527 => "01001010", 16529 => "11000011", 16530 => "11010100", 16531 => "11100000", 16533 => "11001101", 16534 => "11001001", 16538 => "10010001", 16541 => "10011010", 16542 => "01001001", 16543 => "00011010", 16545 => "11010011", 16546 => "00110100", 16548 => "01111110", 16550 => "01111101", 16556 => "00010000", 16557 => "01101011", 16558 => "11011000", 16559 => "01001100", 16560 => "11011001", 16561 => "00111111", 16564 => "01111001", 16565 => "01000101", 16567 => "11100111", 16569 => "11101111", 16570 => "11100010", 16574 => "10110011", 16575 => "10001000", 16579 => "01011011", 16580 => "11111110", 16582 => "10010010", 16583 => "00110111", 16584 => "00001111", 16590 => "01110011", 16594 => "01001001", 16595 => "10111010", 16596 => "00110010", 16597 => "10111100", 16601 => "00101001", 16607 => "11010000", 16612 => "10111001", 16614 => "10000100", 16615 => "00100001", 16617 => "01100110", 16618 => "00100000", 16619 => "10001100", 16620 => "00110011", 16621 => "01001101", 16626 => "11010001", 16627 => "00111111", 16629 => "11011111", 16630 => "11000000", 16632 => "10110000", 16633 => "01100111", 16635 => "01111011", 16636 => "11111101", 16638 => "01011001", 16639 => "10011100", 16640 => "01100100", 16642 => "11010101", 16644 => "11101010", 16647 => "01011000", 16648 => "01111101", 16650 => "00111010", 16651 => "00000011", 16653 => "01010010", 16654 => "00111100", 16656 => "10011001", 16657 => "01011000", 16659 => "00010011", 16661 => "00100001", 16666 => "11101100", 16667 => "01010000", 16669 => "10110101", 16671 => "01110100", 16672 => "11111011", 16673 => "01110101", 16674 => "11111010", 16675 => "01000100", 16676 => "11111100", 16677 => "11100000", 16681 => "01111110", 16683 => "10111001", 16684 => "11011100", 16685 => "11110101", 16690 => "10100000", 16691 => "10101110", 16695 => "11100101", 16697 => "00010101", 16698 => "01001000", 16699 => "10011110", 16703 => "10101111", 16705 => "01100000", 16706 => "01110000", 16707 => "00011001", 16708 => "00111100", 16709 => "01101111", 16711 => "10111000", 16712 => "10101100", 16723 => "00101010", 16724 => "10100000", 16730 => "11100101", 16736 => "01111110", 16738 => "00011111", 16739 => "00011001", 16741 => "10110000", 16745 => "10011011", 16746 => "10111010", 16747 => "01001000", 16749 => "01111010", 16753 => "01001010", 16754 => "11111011", 16755 => "11011101", 16756 => "00001001", 16757 => "11000011", 16758 => "00101100", 16759 => "01001011", 16761 => "01101111", 16763 => "10011010", 16766 => "11100101", 16767 => "01101011", 16769 => "01100100", 16770 => "10110111", 16771 => "10100011", 16774 => "00001011", 16777 => "11101000", 16779 => "00001011", 16780 => "11000001", 16781 => "00011100", 16784 => "01111110", 16789 => "11001101", 16790 => "10010101", 16797 => "11111011", 16800 => "01000110", 16801 => "10011100", 16802 => "01101000", 16804 => "00001110", 16805 => "10011111", 16807 => "10111110", 16809 => "10101000", 16810 => "00111110", 16811 => "10110001", 16814 => "11111111", 16816 => "11101111", 16819 => "01011010", 16822 => "01101110", 16823 => "01001011", 16824 => "10010000", 16826 => "01011110", 16828 => "10010100", 16830 => "11100100", 16831 => "01111110", 16833 => "10001000", 16836 => "00011100", 16838 => "11110111", 16840 => "01110010", 16842 => "01001110", 16846 => "11101001", 16847 => "01100010", 16848 => "11011000", 16849 => "11110111", 16852 => "11111111", 16854 => "01101011", 16855 => "10100110", 16856 => "00011010", 16858 => "00101100", 16859 => "10000111", 16865 => "10010000", 16866 => "11101001", 16869 => "00010110", 16872 => "01001101", 16874 => "10110111", 16875 => "01001001", 16876 => "01100001", 16878 => "11100010", 16880 => "01000100", 16881 => "01011111", 16883 => "11010110", 16884 => "11010001", 16885 => "01010000", 16886 => "11001111", 16889 => "10110111", 16890 => "10011001", 16891 => "11110011", 16894 => "00011101", 16897 => "10100010", 16899 => "11111100", 16901 => "10000000", 16902 => "11111110", 16903 => "11110110", 16909 => "10101100", 16910 => "11010010", 16917 => "10010111", 16919 => "01101111", 16923 => "10000110", 16926 => "11010100", 16933 => "11101001", 16937 => "11001001", 16938 => "10001000", 16942 => "11000010", 16944 => "11100000", 16945 => "11000010", 16947 => "10101011", 16951 => "10101101", 16954 => "10001111", 16955 => "01000110", 16957 => "00101000", 16959 => "00101110", 16962 => "00001010", 16963 => "11100010", 16964 => "01110110", 16965 => "01100000", 16969 => "10010010", 16971 => "00001000", 16974 => "00011111", 16975 => "00110101", 16978 => "11110000", 16980 => "01101100", 16982 => "01000101", 16985 => "00011000", 16987 => "11101010", 16988 => "01000001", 16992 => "01100100", 16994 => "01001011", 16995 => "10111010", 16996 => "11101000", 17001 => "01000001", 17002 => "11011011", 17005 => "00001111", 17006 => "00100000", 17009 => "11001000", 17010 => "00100110", 17011 => "10110100", 17012 => "00011011", 17013 => "11000000", 17014 => "10010111", 17015 => "00010101", 17016 => "00001011", 17020 => "10111111", 17021 => "10101100", 17023 => "01101001", 17024 => "00000100", 17026 => "11111110", 17027 => "01010111", 17028 => "10011110", 17029 => "10111110", 17033 => "01101000", 17036 => "11000011", 17037 => "11100110", 17038 => "11011111", 17040 => "01011101", 17043 => "10010101", 17045 => "01110000", 17048 => "11110001", 17053 => "01101000", 17055 => "11111011", 17057 => "01011111", 17059 => "00000010", 17063 => "10011101", 17066 => "00111100", 17067 => "00100101", 17069 => "11000111", 17072 => "11101101", 17073 => "11111010", 17074 => "01101000", 17075 => "10110010", 17076 => "00010001", 17078 => "01011100", 17080 => "01101001", 17081 => "01001001", 17083 => "00111110", 17084 => "11011001", 17085 => "11110000", 17086 => "11110011", 17088 => "00000100", 17089 => "11010100", 17092 => "00110000", 17093 => "00101001", 17094 => "10100000", 17099 => "10010000", 17100 => "11100010", 17102 => "00000111", 17103 => "10011111", 17105 => "01111010", 17106 => "10010110", 17107 => "10011110", 17109 => "00010011", 17110 => "01001101", 17112 => "01011000", 17117 => "01111100", 17118 => "01000100", 17120 => "00011110", 17121 => "10011100", 17123 => "00111101", 17125 => "01010101", 17127 => "11001110", 17129 => "10000001", 17131 => "11101001", 17134 => "11001111", 17135 => "10001011", 17137 => "10010101", 17139 => "11110000", 17140 => "00011100", 17142 => "11001001", 17143 => "00001001", 17144 => "10101101", 17145 => "00000001", 17147 => "00110010", 17148 => "01101101", 17149 => "10011000", 17150 => "00001000", 17152 => "01010001", 17153 => "10001111", 17155 => "00110100", 17156 => "10110111", 17157 => "00111011", 17160 => "00011000", 17161 => "11011101", 17163 => "10111100", 17164 => "00110111", 17166 => "01011001", 17167 => "10010000", 17168 => "01010010", 17169 => "01110110", 17172 => "11100001", 17174 => "01000101", 17176 => "11011110", 17178 => "00000001", 17179 => "01101111", 17180 => "10111001", 17181 => "01001010", 17182 => "11000100", 17184 => "01100101", 17185 => "10111101", 17186 => "01011010", 17189 => "01000011", 17190 => "10100011", 17192 => "11011111", 17193 => "01010101", 17195 => "01100001", 17199 => "11000011", 17200 => "11111000", 17202 => "10111000", 17207 => "01111011", 17208 => "10101010", 17209 => "01101100", 17210 => "01000110", 17212 => "01110010", 17217 => "00111100", 17218 => "11100000", 17219 => "11111100", 17221 => "01111001", 17227 => "11111001", 17228 => "11111010", 17230 => "00010011", 17232 => "01011001", 17234 => "01000001", 17241 => "11010110", 17245 => "11001110", 17246 => "00111011", 17249 => "01101110", 17250 => "01101100", 17251 => "10110011", 17254 => "01101001", 17255 => "01101000", 17257 => "11000110", 17259 => "11110000", 17265 => "10110110", 17266 => "00000100", 17268 => "11011010", 17270 => "10101001", 17271 => "10110011", 17272 => "00011110", 17276 => "11100110", 17277 => "11111100", 17279 => "10110101", 17281 => "11010011", 17283 => "10011010", 17286 => "11011010", 17287 => "10110001", 17289 => "10111011", 17291 => "11010010", 17293 => "11100010", 17295 => "01010000", 17296 => "00010101", 17299 => "01111100", 17302 => "00110110", 17304 => "10101001", 17305 => "10101101", 17306 => "01110110", 17308 => "00000001", 17310 => "00010010", 17312 => "00101110", 17313 => "10001111", 17314 => "00000010", 17316 => "11100011", 17318 => "00111110", 17323 => "01100110", 17324 => "00101001", 17326 => "01111111", 17330 => "10000100", 17331 => "00000001", 17332 => "10001110", 17333 => "00000001", 17334 => "01010101", 17335 => "10110101", 17336 => "00100000", 17337 => "00111000", 17338 => "01110000", 17339 => "10011111", 17341 => "00100000", 17342 => "10001000", 17345 => "11000001", 17346 => "11001111", 17348 => "01111100", 17351 => "11000101", 17352 => "11010101", 17353 => "10000100", 17355 => "10111110", 17356 => "11001001", 17357 => "11001100", 17358 => "11110111", 17359 => "11010111", 17360 => "01000110", 17361 => "11001010", 17365 => "10001001", 17366 => "00111100", 17368 => "01000110", 17370 => "01111110", 17371 => "11101101", 17372 => "10100001", 17373 => "00101100", 17375 => "00101011", 17379 => "00101100", 17380 => "00110000", 17381 => "00001111", 17382 => "10001101", 17383 => "01111101", 17387 => "01001110", 17388 => "01110001", 17390 => "11111001", 17392 => "00111100", 17393 => "01101011", 17394 => "01000101", 17396 => "11010011", 17397 => "00000001", 17399 => "10111111", 17400 => "10101000", 17402 => "01010111", 17403 => "11010111", 17404 => "10111000", 17410 => "11000110", 17416 => "00101010", 17421 => "11111011", 17422 => "11110011", 17423 => "00001000", 17430 => "11111000", 17432 => "00010110", 17435 => "10011011", 17436 => "10110111", 17437 => "10110001", 17438 => "00010000", 17443 => "11101010", 17444 => "10111000", 17445 => "11000110", 17446 => "10010111", 17450 => "00000111", 17452 => "00001100", 17455 => "00011000", 17458 => "10000100", 17459 => "00011011", 17461 => "10000111", 17463 => "10001010", 17467 => "01100010", 17468 => "11101011", 17469 => "01101000", 17472 => "01010000", 17473 => "10100010", 17474 => "11000110", 17475 => "01100011", 17478 => "10010001", 17481 => "11011111", 17483 => "10111111", 17485 => "00000100", 17488 => "10110111", 17489 => "00010001", 17493 => "10010000", 17494 => "01100000", 17495 => "00001101", 17499 => "11001110", 17501 => "10110100", 17502 => "10001101", 17503 => "01001111", 17504 => "01110101", 17505 => "00011111", 17509 => "11000000", 17511 => "01010000", 17512 => "01101001", 17513 => "11000101", 17514 => "10101000", 17515 => "00111011", 17516 => "00101000", 17518 => "01001010", 17520 => "00110011", 17521 => "00000110", 17522 => "10001101", 17523 => "01001110", 17524 => "10000110", 17525 => "00111010", 17526 => "00100010", 17527 => "11101111", 17530 => "01100010", 17534 => "00110100", 17537 => "10111011", 17538 => "00100011", 17539 => "01101110", 17541 => "00101111", 17542 => "11000000", 17545 => "10101111", 17546 => "00111000", 17548 => "11011100", 17550 => "11000000", 17551 => "10001111", 17556 => "10001100", 17559 => "01011000", 17561 => "11100011", 17563 => "00010100", 17564 => "11000000", 17565 => "00111101", 17566 => "00100011", 17567 => "00100110", 17569 => "01010011", 17574 => "10101010", 17575 => "11110001", 17577 => "00010101", 17579 => "00100100", 17580 => "01110110", 17585 => "00100000", 17587 => "11000000", 17588 => "00000010", 17589 => "01100010", 17590 => "00101101", 17591 => "11110100", 17592 => "00001001", 17593 => "10111001", 17594 => "10011100", 17595 => "00010011", 17596 => "11011110", 17600 => "01101100", 17603 => "00110000", 17604 => "10010001", 17605 => "01101001", 17606 => "10011111", 17609 => "10101011", 17612 => "01101011", 17613 => "01010010", 17615 => "10100000", 17616 => "11000101", 17617 => "11110111", 17618 => "10101011", 17621 => "01100100", 17623 => "01111101", 17624 => "01000100", 17629 => "11000001", 17630 => "11101011", 17631 => "01000110", 17633 => "01101011", 17639 => "01010000", 17640 => "10101010", 17641 => "00110111", 17642 => "11101101", 17643 => "10101010", 17644 => "10001001", 17645 => "01100011", 17647 => "11100010", 17650 => "10111101", 17651 => "10101110", 17656 => "01110010", 17657 => "00010011", 17659 => "11110110", 17662 => "00100001", 17663 => "00011010", 17664 => "10010111", 17667 => "01010010", 17669 => "01111111", 17671 => "11011001", 17672 => "00001000", 17674 => "00100101", 17677 => "10101010", 17680 => "00011011", 17681 => "01110100", 17682 => "00011010", 17685 => "01010001", 17688 => "00111110", 17690 => "00011100", 17692 => "01100111", 17693 => "11011110", 17695 => "11101010", 17696 => "00101101", 17701 => "11111111", 17702 => "00111010", 17708 => "01001111", 17711 => "01001011", 17713 => "01101110", 17714 => "01000111", 17720 => "11110001", 17721 => "00000110", 17722 => "01100111", 17724 => "00111111", 17725 => "01011100", 17732 => "00101011", 17735 => "00111010", 17737 => "01111100", 17741 => "00011100", 17743 => "10001110", 17744 => "01010101", 17745 => "01010011", 17747 => "00111111", 17748 => "01100111", 17751 => "10011100", 17752 => "00011000", 17753 => "11101011", 17754 => "11000111", 17758 => "00110000", 17760 => "10101111", 17768 => "11011101", 17769 => "11101111", 17770 => "00101100", 17771 => "00011111", 17772 => "10001011", 17774 => "01110111", 17776 => "11001010", 17778 => "10000010", 17779 => "00001001", 17782 => "11101000", 17783 => "00110101", 17785 => "10010110", 17786 => "10000011", 17787 => "11101111", 17788 => "00011100", 17790 => "01011010", 17791 => "11011100", 17792 => "10000000", 17796 => "10010001", 17797 => "00010000", 17798 => "00110110", 17799 => "01000111", 17800 => "00001111", 17801 => "01100110", 17803 => "10100010", 17809 => "11111110", 17810 => "01100110", 17812 => "01010011", 17813 => "10101010", 17815 => "01110010", 17816 => "11100010", 17817 => "10010101", 17819 => "11000101", 17820 => "11100011", 17822 => "00100101", 17823 => "11111000", 17825 => "01001110", 17826 => "11111001", 17829 => "01001010", 17831 => "11000000", 17834 => "01110100", 17836 => "10010000", 17837 => "11100001", 17839 => "10100110", 17849 => "01111111", 17850 => "11101111", 17853 => "00100001", 17855 => "00111101", 17856 => "00010100", 17858 => "11000001", 17859 => "01111101", 17860 => "01111000", 17861 => "11011111", 17862 => "01100001", 17863 => "01101001", 17864 => "00100100", 17867 => "11101100", 17870 => "01000011", 17871 => "00011111", 17873 => "11010011", 17876 => "00101011", 17877 => "11100000", 17878 => "00110001", 17881 => "10000101", 17882 => "10010110", 17885 => "11101101", 17889 => "11010001", 17890 => "01010010", 17891 => "11111001", 17894 => "10001110", 17895 => "11111000", 17896 => "11010000", 17897 => "10101010", 17901 => "10000111", 17902 => "10111011", 17903 => "11000011", 17905 => "10110011", 17907 => "00000011", 17911 => "11010100", 17912 => "00100100", 17913 => "01100100", 17914 => "11010100", 17915 => "01011111", 17916 => "01010111", 17917 => "11111010", 17919 => "01111001", 17920 => "11101100", 17921 => "01000100", 17923 => "11111110", 17926 => "10110110", 17927 => "00110110", 17928 => "10000011", 17929 => "11110001", 17930 => "11000000", 17932 => "00111111", 17933 => "11000101", 17934 => "10001011", 17936 => "00010101", 17938 => "00010101", 17943 => "10101100", 17948 => "00011011", 17949 => "00110100", 17950 => "00100010", 17951 => "00101000", 17952 => "10110001", 17953 => "01100110", 17954 => "00011111", 17955 => "01011001", 17956 => "00101001", 17962 => "10011111", 17965 => "11001010", 17966 => "00111110", 17973 => "00101110", 17974 => "01001000", 17975 => "11110011", 17976 => "01000111", 17978 => "00001001", 17979 => "00011000", 17982 => "10011000", 17983 => "11000001", 17985 => "01100101", 17988 => "00111100", 17989 => "00011101", 17990 => "00100110", 17993 => "00010010", 17994 => "10011110", 17995 => "11100000", 17998 => "11001010", 17999 => "00100011", 18000 => "10000101", 18001 => "10100011", 18002 => "11100100", 18003 => "11011111", 18005 => "00001110", 18008 => "00101110", 18009 => "10101011", 18012 => "01110110", 18015 => "00011001", 18019 => "11100010", 18028 => "10000000", 18029 => "11100101", 18032 => "11110110", 18034 => "01001101", 18036 => "11001101", 18037 => "01010110", 18038 => "11001100", 18039 => "11010011", 18042 => "01100110", 18045 => "01101001", 18049 => "10001001", 18052 => "00000100", 18053 => "00110001", 18054 => "01000101", 18056 => "10100000", 18057 => "10111110", 18058 => "11011011", 18060 => "11111111", 18062 => "01100001", 18063 => "01011001", 18064 => "01100011", 18068 => "11000000", 18070 => "11110100", 18072 => "01101110", 18073 => "11110100", 18074 => "10101100", 18075 => "00101110", 18077 => "10010100", 18081 => "10010011", 18082 => "10000110", 18083 => "01100011", 18090 => "11101100", 18091 => "11001011", 18093 => "11011011", 18094 => "11000100", 18097 => "11010100", 18098 => "10110001", 18100 => "00010001", 18101 => "11100111", 18103 => "01110111", 18104 => "11011011", 18105 => "01100011", 18107 => "01110111", 18110 => "11100010", 18112 => "01001111", 18114 => "01011111", 18115 => "00010110", 18116 => "10100110", 18117 => "01010110", 18118 => "00000101", 18119 => "10110110", 18121 => "11000110", 18124 => "10111111", 18126 => "00101011", 18127 => "10101101", 18128 => "10010100", 18129 => "10111001", 18131 => "01110101", 18132 => "11001000", 18133 => "01100100", 18134 => "01110101", 18137 => "00010011", 18138 => "00101001", 18139 => "01000011", 18141 => "10110011", 18144 => "00010100", 18147 => "00000100", 18149 => "11101010", 18150 => "11111100", 18153 => "10100101", 18154 => "11111100", 18155 => "10000010", 18157 => "01111001", 18159 => "01110000", 18160 => "00110111", 18162 => "00011110", 18163 => "01010111", 18164 => "01100101", 18168 => "10011110", 18169 => "10001101", 18172 => "10010100", 18180 => "01100010", 18182 => "10101000", 18183 => "11000001", 18187 => "00111010", 18188 => "00100001", 18189 => "11110110", 18191 => "00100010", 18194 => "00011111", 18199 => "11100000", 18200 => "10100011", 18201 => "10100111", 18202 => "00000011", 18204 => "10100101", 18211 => "11111000", 18213 => "00110101", 18214 => "11111101", 18215 => "00011100", 18216 => "01010000", 18218 => "10010010", 18223 => "00101110", 18224 => "10111111", 18226 => "10011110", 18231 => "00000001", 18232 => "00100000", 18234 => "10100101", 18235 => "01111010", 18238 => "11101101", 18239 => "11111011", 18245 => "00010101", 18247 => "00100010", 18249 => "11010110", 18251 => "10111110", 18255 => "01011111", 18257 => "00010110", 18258 => "00110110", 18261 => "10110001", 18262 => "00010011", 18265 => "00100010", 18266 => "01101100", 18268 => "00000110", 18269 => "11100110", 18270 => "01001000", 18272 => "01111101", 18273 => "11001010", 18276 => "00011101", 18277 => "11001101", 18280 => "01000100", 18282 => "01011111", 18287 => "11111011", 18288 => "11001101", 18290 => "01111010", 18292 => "10101100", 18295 => "11100000", 18297 => "10101110", 18300 => "11011101", 18301 => "00011101", 18302 => "10110000", 18304 => "11001000", 18306 => "10010010", 18308 => "00001100", 18309 => "00110011", 18312 => "01000111", 18313 => "11111111", 18316 => "01011001", 18318 => "11011011", 18319 => "00011010", 18321 => "10011000", 18325 => "00100111", 18326 => "10110110", 18328 => "11101110", 18329 => "10101011", 18330 => "10001010", 18331 => "11011101", 18334 => "11000110", 18338 => "01001101", 18339 => "00000100", 18340 => "11010100", 18344 => "00011011", 18345 => "01111011", 18348 => "01011101", 18355 => "01110100", 18357 => "10010100", 18358 => "10010001", 18359 => "01111000", 18361 => "11100111", 18363 => "01101100", 18365 => "01111011", 18369 => "00100000", 18371 => "10000011", 18372 => "10011010", 18373 => "11101011", 18374 => "11100001", 18377 => "10111111", 18385 => "01111100", 18386 => "11011111", 18389 => "11110001", 18393 => "11000111", 18394 => "11110110", 18395 => "01111011", 18396 => "00100010", 18397 => "01100010", 18398 => "10100111", 18399 => "00001011", 18400 => "01100111", 18402 => "00010010", 18404 => "00011100", 18405 => "00100100", 18406 => "10111010", 18407 => "10000000", 18409 => "01000011", 18411 => "10010000", 18412 => "01101000", 18413 => "01100100", 18414 => "10111110", 18418 => "10010100", 18419 => "11011010", 18421 => "11111011", 18423 => "11111010", 18425 => "11110110", 18426 => "00101000", 18428 => "00010111", 18430 => "11101010", 18434 => "10101010", 18435 => "01101000", 18436 => "01010100", 18443 => "11000011", 18445 => "00001010", 18448 => "11011101", 18449 => "11001111", 18451 => "10110111", 18452 => "10000000", 18453 => "11100000", 18454 => "01010000", 18455 => "11101111", 18458 => "01000111", 18464 => "01101111", 18467 => "01000011", 18469 => "01111111", 18471 => "11010100", 18472 => "11111101", 18473 => "01100111", 18477 => "00011100", 18480 => "00110101", 18481 => "10001000", 18482 => "01100111", 18487 => "01101101", 18488 => "10011110", 18490 => "00001110", 18491 => "00111100", 18494 => "10101000", 18495 => "10100010", 18496 => "11000001", 18499 => "01000001", 18501 => "11010000", 18502 => "10011100", 18503 => "11011111", 18505 => "00011011", 18506 => "11011011", 18507 => "11000010", 18509 => "00011100", 18510 => "01001000", 18511 => "00111101", 18512 => "10101111", 18515 => "10010111", 18516 => "10001100", 18517 => "10001001", 18518 => "11010011", 18520 => "01001000", 18522 => "00110101", 18523 => "00111001", 18525 => "00000100", 18526 => "11000001", 18528 => "11010001", 18529 => "10000010", 18538 => "01010101", 18539 => "01001111", 18540 => "11011110", 18541 => "11110100", 18542 => "01110001", 18543 => "01110010", 18544 => "10101001", 18546 => "10001001", 18547 => "11110101", 18550 => "11111101", 18551 => "10111011", 18552 => "00111001", 18557 => "11101001", 18558 => "11111110", 18559 => "00001111", 18560 => "11110100", 18564 => "01010101", 18565 => "01001110", 18567 => "11000110", 18568 => "10011000", 18572 => "10000101", 18575 => "11100011", 18577 => "01100111", 18579 => "11011010", 18581 => "00100100", 18582 => "01001001", 18583 => "00011000", 18584 => "01010100", 18585 => "11001101", 18586 => "10110100", 18588 => "11111111", 18590 => "10110011", 18591 => "11000010", 18592 => "00011001", 18594 => "00100011", 18597 => "01011100", 18602 => "10001010", 18604 => "01101011", 18605 => "11100111", 18607 => "00110101", 18609 => "00010000", 18612 => "11101011", 18614 => "01111010", 18615 => "10010010", 18617 => "01110010", 18618 => "11011011", 18623 => "01110000", 18624 => "11001110", 18627 => "10101011", 18628 => "01101001", 18631 => "10110110", 18634 => "01111011", 18635 => "00001101", 18636 => "00011100", 18638 => "01010110", 18639 => "11000101", 18640 => "10001011", 18641 => "11110111", 18642 => "10000000", 18645 => "11100010", 18647 => "01001010", 18649 => "10100010", 18650 => "10100000", 18652 => "01111010", 18656 => "00101000", 18658 => "11111010", 18659 => "11100101", 18661 => "10000011", 18663 => "10011110", 18667 => "10001000", 18668 => "11001111", 18669 => "00010111", 18670 => "11011110", 18671 => "00111100", 18672 => "10010011", 18673 => "11111110", 18674 => "01011111", 18681 => "01001010", 18682 => "00010000", 18685 => "01111010", 18686 => "10110000", 18687 => "10001011", 18688 => "01100101", 18692 => "11100100", 18698 => "01101100", 18699 => "11000000", 18701 => "11110000", 18702 => "00000100", 18703 => "10001011", 18705 => "10001010", 18709 => "10100000", 18711 => "10000000", 18712 => "11001100", 18713 => "01010111", 18714 => "11000000", 18715 => "00111010", 18716 => "11100001", 18719 => "01010110", 18720 => "10110000", 18721 => "11001001", 18722 => "01001100", 18725 => "01011100", 18726 => "01110011", 18729 => "01110110", 18732 => "00010110", 18734 => "00001101", 18745 => "10011001", 18748 => "00010010", 18749 => "10001000", 18750 => "11000001", 18751 => "11010110", 18754 => "10001001", 18755 => "11111100", 18756 => "00110001", 18757 => "01011000", 18758 => "11101011", 18760 => "01100011", 18766 => "11010100", 18768 => "11001000", 18769 => "01110100", 18770 => "01111011", 18776 => "10011101", 18780 => "01011000", 18784 => "11010100", 18785 => "00011110", 18787 => "11011110", 18788 => "00011000", 18794 => "11100111", 18797 => "00101000", 18801 => "11111000", 18802 => "10001000", 18806 => "10010111", 18809 => "11010000", 18812 => "01101001", 18813 => "11011101", 18814 => "01011010", 18820 => "00110100", 18821 => "01110100", 18823 => "10000111", 18824 => "00101101", 18829 => "10100101", 18830 => "11010001", 18832 => "11101011", 18835 => "01101001", 18838 => "00101010", 18839 => "01000100", 18840 => "10000001", 18843 => "11010001", 18844 => "11010110", 18845 => "10011011", 18850 => "01010100", 18851 => "00011111", 18852 => "00010101", 18853 => "01011000", 18856 => "11000010", 18859 => "10111100", 18860 => "01100110", 18862 => "11101001", 18866 => "11010111", 18868 => "01010111", 18869 => "11101100", 18873 => "00001001", 18874 => "10011011", 18875 => "01011100", 18876 => "10101111", 18880 => "01000101", 18883 => "11100000", 18885 => "10100101", 18887 => "00100110", 18889 => "01001111", 18894 => "10111000", 18895 => "00110111", 18899 => "01010100", 18900 => "10010110", 18905 => "01111010", 18907 => "01010010", 18909 => "01110110", 18910 => "00100000", 18911 => "01100001", 18912 => "00111000", 18913 => "00110111", 18915 => "11110001", 18916 => "10110101", 18922 => "01101101", 18923 => "11010001", 18926 => "01111011", 18928 => "01100101", 18931 => "00111010", 18935 => "00010100", 18936 => "00111111", 18938 => "01000111", 18941 => "10001010", 18942 => "00011010", 18944 => "11100101", 18945 => "00011111", 18947 => "11011101", 18948 => "01110001", 18949 => "10010001", 18953 => "01010001", 18955 => "01011011", 18960 => "10111110", 18961 => "10100100", 18963 => "11010101", 18964 => "01111111", 18965 => "00001110", 18967 => "00100000", 18970 => "00010000", 18971 => "01111011", 18975 => "01111110", 18976 => "11011011", 18981 => "00110011", 18982 => "01111001", 18983 => "01111011", 18984 => "11000100", 18988 => "01000101", 18992 => "10011101", 18993 => "10000010", 18995 => "00111000", 18998 => "11010000", 19001 => "01111100", 19003 => "01010110", 19005 => "01110011", 19006 => "10011101", 19010 => "10000100", 19011 => "10111100", 19017 => "10001101", 19018 => "01111100", 19019 => "01010101", 19020 => "00100001", 19022 => "01001101", 19023 => "01001111", 19025 => "10010110", 19027 => "01000100", 19028 => "10100010", 19029 => "00110101", 19034 => "00110100", 19035 => "11000110", 19036 => "10011011", 19037 => "10000011", 19040 => "00100011", 19041 => "11011110", 19042 => "00110110", 19043 => "00110010", 19045 => "01010000", 19046 => "10000101", 19048 => "00010010", 19050 => "01001100", 19051 => "01010110", 19053 => "01011101", 19054 => "01101001", 19055 => "00111100", 19057 => "01100101", 19060 => "00011000", 19061 => "01000101", 19062 => "10111110", 19066 => "11100110", 19067 => "01110011", 19069 => "01010100", 19071 => "10110101", 19072 => "11011100", 19074 => "11001001", 19081 => "00000111", 19082 => "10111000", 19084 => "00100011", 19087 => "11000100", 19089 => "10110000", 19090 => "11100000", 19091 => "10010001", 19093 => "10000111", 19096 => "11100110", 19098 => "11110111", 19100 => "00001100", 19103 => "11100001", 19106 => "00001000", 19109 => "11000111", 19110 => "11000010", 19113 => "01011001", 19115 => "10000010", 19118 => "00101110", 19119 => "11100001", 19120 => "01010010", 19124 => "00111100", 19126 => "01101110", 19129 => "01101101", 19134 => "01101010", 19136 => "00101101", 19140 => "10011101", 19141 => "11001100", 19146 => "01111010", 19147 => "00010000", 19156 => "00100010", 19158 => "01101001", 19159 => "11100000", 19164 => "01110001", 19166 => "10010110", 19167 => "11001101", 19168 => "01110101", 19173 => "10001010", 19177 => "01100110", 19179 => "10001001", 19181 => "00001111", 19182 => "01100000", 19190 => "11111001", 19191 => "11101010", 19193 => "00011110", 19195 => "10011100", 19196 => "10100110", 19197 => "00110111", 19199 => "10100010", 19200 => "10010110", 19202 => "10110101", 19203 => "11101100", 19204 => "10000011", 19205 => "00100010", 19207 => "11010111", 19208 => "11111001", 19209 => "11000010", 19217 => "10011010", 19220 => "01011110", 19222 => "11100000", 19223 => "00110001", 19226 => "10111101", 19231 => "01000101", 19233 => "00110011", 19234 => "11001111", 19236 => "01010100", 19238 => "00000111", 19239 => "11111101", 19242 => "00010001", 19243 => "01110011", 19244 => "01111100", 19246 => "11001011", 19247 => "00001100", 19248 => "11001000", 19250 => "10011010", 19253 => "01000000", 19254 => "10111110", 19256 => "10000111", 19257 => "10010101", 19259 => "01011100", 19262 => "00110110", 19263 => "01110110", 19266 => "11010011", 19268 => "11000010", 19269 => "01110001", 19270 => "11101011", 19271 => "10110011", 19272 => "00010001", 19273 => "01001111", 19275 => "01100111", 19280 => "11011010", 19282 => "00000001", 19283 => "00100101", 19284 => "01111011", 19285 => "01110010", 19286 => "00100100", 19288 => "00010101", 19290 => "01111010", 19291 => "00010000", 19295 => "11111100", 19296 => "00110000", 19297 => "10101000", 19298 => "11100100", 19300 => "00110000", 19301 => "00011111", 19304 => "01100100", 19306 => "11101111", 19307 => "11001001", 19308 => "00100101", 19309 => "10011001", 19310 => "11100000", 19319 => "10010100", 19320 => "01110110", 19322 => "00001001", 19324 => "11101100", 19326 => "11001100", 19329 => "11001111", 19337 => "00100010", 19345 => "01110111", 19349 => "00010101", 19351 => "00011110", 19356 => "11000000", 19357 => "01010001", 19363 => "01110000", 19365 => "11101100", 19370 => "00011000", 19371 => "00011110", 19372 => "10101000", 19373 => "11010010", 19374 => "10010001", 19375 => "01101001", 19376 => "00101100", 19377 => "10001110", 19378 => "10101001", 19379 => "10000110", 19381 => "11000111", 19383 => "00111010", 19386 => "10011001", 19389 => "01111011", 19391 => "00001010", 19392 => "10100101", 19397 => "10111001", 19398 => "11000001", 19400 => "11110001", 19401 => "11111010", 19402 => "00001000", 19404 => "01001001", 19406 => "11000100", 19407 => "00111000", 19408 => "10111101", 19410 => "11111100", 19411 => "10010100", 19416 => "11011010", 19417 => "01010000", 19418 => "01100000", 19419 => "00000011", 19420 => "10011111", 19421 => "11101101", 19422 => "01110100", 19424 => "10010101", 19425 => "01001001", 19427 => "00000100", 19428 => "00100101", 19434 => "00101010", 19442 => "00100001", 19443 => "01101011", 19445 => "11110001", 19446 => "11001100", 19448 => "10111000", 19450 => "00001101", 19451 => "00011000", 19456 => "00011010", 19460 => "01111101", 19462 => "10110111", 19465 => "10100001", 19466 => "10110111", 19470 => "10110111", 19473 => "10010101", 19474 => "10110010", 19475 => "01000100", 19478 => "10111101", 19479 => "11001111", 19481 => "01001110", 19482 => "10101011", 19483 => "00001010", 19484 => "10100101", 19487 => "10000111", 19488 => "01010111", 19489 => "11010101", 19491 => "11100011", 19494 => "00100100", 19497 => "00000011", 19500 => "00100110", 19501 => "11011111", 19502 => "10000011", 19503 => "00001010", 19506 => "10100110", 19508 => "00100001", 19510 => "00000100", 19511 => "10010001", 19514 => "11001110", 19516 => "00011101", 19517 => "01101011", 19519 => "00110000", 19521 => "10110100", 19522 => "01000011", 19524 => "00001001", 19526 => "11101110", 19528 => "01110010", 19529 => "10011101", 19531 => "01110010", 19532 => "10110011", 19535 => "01000001", 19536 => "00010000", 19540 => "11111110", 19541 => "01110011", 19542 => "01010000", 19543 => "10111000", 19544 => "10101110", 19545 => "11110110", 19546 => "10010001", 19549 => "00001000", 19550 => "01100101", 19551 => "10101110", 19553 => "00011010", 19554 => "11000000", 19556 => "10001011", 19557 => "01101001", 19562 => "11001110", 19563 => "11111011", 19564 => "11100000", 19568 => "10100010", 19570 => "00001010", 19572 => "11011001", 19573 => "00011110", 19574 => "10010010", 19575 => "10011101", 19579 => "00111000", 19580 => "10110010", 19581 => "10000000", 19583 => "01001001", 19584 => "01101001", 19586 => "10111111", 19587 => "11101011", 19589 => "10010010", 19590 => "11001011", 19591 => "11010101", 19592 => "00100111", 19593 => "00101100", 19595 => "11110010", 19596 => "11110111", 19600 => "00010100", 19602 => "01100011", 19605 => "00111110", 19613 => "00001101", 19614 => "11001001", 19617 => "01101011", 19619 => "01100011", 19620 => "11001011", 19621 => "10001110", 19622 => "10101010", 19623 => "00010100", 19626 => "00001001", 19628 => "11010111", 19630 => "00100101", 19633 => "00100101", 19634 => "01010101", 19638 => "10010001", 19643 => "11001010", 19645 => "01111101", 19647 => "00100001", 19649 => "10111100", 19650 => "01101000", 19651 => "11000001", 19653 => "01110001", 19655 => "11000010", 19658 => "01111101", 19661 => "01100000", 19663 => "10100011", 19669 => "11100110", 19670 => "11000011", 19672 => "11011000", 19673 => "10111000", 19674 => "11010100", 19675 => "00101111", 19676 => "00111000", 19677 => "11001111", 19678 => "11100100", 19679 => "10000100", 19682 => "01111010", 19691 => "10001111", 19693 => "00011000", 19697 => "11010100", 19698 => "10101110", 19699 => "01110101", 19700 => "10111100", 19701 => "10001001", 19702 => "01100101", 19703 => "01011010", 19707 => "10110000", 19709 => "11111110", 19710 => "01100011", 19713 => "10101001", 19715 => "00010100", 19716 => "00010110", 19718 => "11100000", 19720 => "11011000", 19723 => "00100110", 19727 => "01010101", 19736 => "01000010", 19743 => "10101010", 19744 => "01001101", 19745 => "01010100", 19746 => "00110110", 19748 => "10101000", 19749 => "01100101", 19753 => "10110011", 19754 => "00101111", 19755 => "01010101", 19761 => "01101010", 19762 => "11010010", 19763 => "10100100", 19764 => "11011101", 19766 => "10011110", 19767 => "11101001", 19770 => "01110000", 19772 => "00000110", 19773 => "10110010", 19774 => "11011010", 19775 => "01101100", 19776 => "00010111", 19777 => "11011010", 19778 => "11000110", 19781 => "11111110", 19784 => "11100000", 19785 => "00101100", 19786 => "00100000", 19788 => "01101101", 19790 => "01010010", 19791 => "01100000", 19792 => "00011100", 19793 => "11110011", 19795 => "11111101", 19796 => "10111000", 19797 => "10101001", 19798 => "10101110", 19801 => "00100111", 19802 => "11001101", 19804 => "00100111", 19805 => "00100100", 19806 => "10100010", 19810 => "10111111", 19811 => "11000001", 19813 => "00010101", 19814 => "01010100", 19815 => "01100010", 19816 => "01110011", 19825 => "01000100", 19827 => "11101000", 19828 => "01101000", 19830 => "11110101", 19832 => "01100111", 19835 => "10011011", 19838 => "11000001", 19843 => "11001011", 19845 => "11101101", 19847 => "11011011", 19849 => "01001011", 19850 => "11011010", 19851 => "11111010", 19853 => "01001111", 19855 => "01010100", 19856 => "01110111", 19857 => "10000100", 19859 => "10011001", 19860 => "10110011", 19862 => "01000000", 19864 => "10110101", 19867 => "10010001", 19868 => "10101011", 19872 => "00011011", 19876 => "11000100", 19877 => "11000001", 19878 => "00100001", 19879 => "10010001", 19881 => "01010100", 19882 => "01001100", 19883 => "01010011", 19885 => "11110000", 19886 => "10110011", 19888 => "01110001", 19889 => "00000001", 19890 => "10100011", 19891 => "10000010", 19892 => "11001000", 19893 => "10111010", 19895 => "00110100", 19898 => "11011110", 19901 => "10110010", 19902 => "00111010", 19903 => "11100011", 19908 => "11011111", 19910 => "00001011", 19914 => "10000000", 19916 => "11000011", 19917 => "01000101", 19918 => "00010111", 19921 => "01111100", 19925 => "01100111", 19926 => "10101100", 19927 => "01101011", 19931 => "00011010", 19935 => "10011111", 19938 => "11111101", 19939 => "01010001", 19942 => "11111101", 19943 => "11100011", 19946 => "01000010", 19950 => "11001000", 19951 => "11100111", 19952 => "01101110", 19953 => "01101001", 19954 => "00001100", 19956 => "10010011", 19957 => "10011000", 19959 => "10110010", 19960 => "00111111", 19961 => "01110010", 19968 => "10100100", 19970 => "01011010", 19971 => "10011100", 19973 => "11001011", 19974 => "10101111", 19975 => "01110101", 19976 => "01100100", 19977 => "01011010", 19979 => "10001010", 19980 => "01000111", 19981 => "00101101", 19984 => "00001001", 19985 => "10001101", 19987 => "00010110", 19988 => "10000110", 19989 => "00010011", 19990 => "10110001", 19995 => "01001011", 19996 => "00101101", 19997 => "11010101", 20000 => "00000100", 20001 => "00100010", 20002 => "10101100", 20004 => "00000111", 20006 => "00101110", 20009 => "10001000", 20010 => "00100010", 20011 => "01100101", 20013 => "11111001", 20019 => "01011111", 20023 => "11110100", 20027 => "11111110", 20029 => "11001100", 20030 => "11100110", 20032 => "01000010", 20036 => "11111011", 20037 => "01000011", 20039 => "11100110", 20043 => "10011111", 20044 => "01011010", 20047 => "00001110", 20057 => "00100011", 20059 => "10101100", 20060 => "10001111", 20062 => "10011000", 20064 => "10000010", 20065 => "10110010", 20068 => "11101001", 20070 => "01100110", 20071 => "00111010", 20074 => "01010010", 20076 => "00110000", 20077 => "10010010", 20081 => "00010110", 20084 => "10100110", 20086 => "00011101", 20087 => "01011001", 20088 => "01100101", 20089 => "10001100", 20090 => "00001001", 20091 => "11001111", 20095 => "10110110", 20096 => "11110010", 20097 => "00101001", 20101 => "10101111", 20102 => "11101111", 20104 => "00101010", 20105 => "11111101", 20108 => "00000011", 20110 => "00010101", 20111 => "00100111", 20112 => "01110110", 20114 => "11010100", 20117 => "11011110", 20121 => "01110101", 20124 => "10110000", 20125 => "00111110", 20128 => "00100000", 20130 => "10110001", 20131 => "10001010", 20134 => "11110000", 20136 => "11111110", 20137 => "01001101", 20138 => "11111111", 20141 => "00100100", 20142 => "10101010", 20145 => "10110001", 20148 => "11101101", 20150 => "01110110", 20151 => "11001110", 20153 => "00110010", 20155 => "10101100", 20156 => "00100101", 20157 => "01010010", 20164 => "01110101", 20165 => "00000010", 20166 => "01101001", 20168 => "11011011", 20169 => "00001000", 20170 => "11110100", 20172 => "11001111", 20174 => "00001101", 20175 => "01010010", 20183 => "01001111", 20185 => "11111111", 20188 => "01011000", 20189 => "10010110", 20190 => "01011010", 20191 => "10000001", 20192 => "11100110", 20193 => "10111101", 20195 => "10010111", 20198 => "10100110", 20200 => "01100100", 20203 => "00110000", 20204 => "10011111", 20206 => "11000000", 20207 => "11000010", 20210 => "00011100", 20213 => "11110000", 20214 => "10110001", 20216 => "01010001", 20218 => "11001000", 20219 => "11011000", 20220 => "01110100", 20224 => "00011010", 20225 => "10000000", 20230 => "00101011", 20235 => "11000011", 20237 => "11101001", 20238 => "00111000", 20249 => "10011100", 20251 => "11110001", 20252 => "11001111", 20253 => "11011001", 20256 => "11001101", 20259 => "10110011", 20264 => "10010000", 20266 => "10010010", 20267 => "00001011", 20268 => "11100100", 20270 => "01101100", 20272 => "10001100", 20273 => "10111100", 20274 => "10101100", 20276 => "10111011", 20279 => "10001110", 20280 => "10111000", 20282 => "10110101", 20283 => "10001010", 20284 => "10110111", 20285 => "10001001", 20286 => "00010100", 20288 => "00100011", 20292 => "11100001", 20294 => "10100101", 20299 => "01101110", 20300 => "00100100", 20304 => "00010110", 20306 => "10010100", 20307 => "10011110", 20311 => "10110100", 20315 => "01111100", 20316 => "11000101", 20317 => "11001110", 20321 => "00010100", 20322 => "00010110", 20324 => "10111011", 20328 => "01000001", 20329 => "01111000", 20330 => "00111111", 20334 => "00001010", 20337 => "11010000", 20338 => "00011101", 20343 => "00010010", 20344 => "00111000", 20345 => "10000100", 20347 => "11000110", 20349 => "00001011", 20350 => "01011110", 20351 => "00100011", 20353 => "11100010", 20354 => "01101100", 20356 => "00001111", 20359 => "10001011", 20361 => "00111010", 20363 => "01100011", 20364 => "10000011", 20369 => "00110110", 20374 => "11001001", 20375 => "10110111", 20377 => "00111100", 20378 => "11111110", 20379 => "01001010", 20382 => "00010110", 20383 => "10110000", 20386 => "00001101", 20387 => "11101010", 20388 => "00001100", 20391 => "11110110", 20394 => "00110100", 20398 => "01010010", 20399 => "00000001", 20403 => "00110101", 20405 => "01010001", 20406 => "11000001", 20407 => "11001000", 20409 => "00001000", 20410 => "01100111", 20411 => "00011000", 20413 => "00101110", 20414 => "01001000", 20415 => "11110100", 20417 => "11111100", 20419 => "00011110", 20422 => "00110001", 20425 => "10111010", 20426 => "00111010", 20428 => "01010101", 20429 => "11000110", 20433 => "01000011", 20434 => "01000000", 20436 => "10001111", 20439 => "01100001", 20441 => "00100111", 20442 => "00101101", 20446 => "01011011", 20448 => "01010011", 20449 => "11011101", 20450 => "01010111", 20451 => "10011101", 20452 => "11110101", 20455 => "01110101", 20456 => "00001011", 20458 => "10110010", 20459 => "01110011", 20462 => "01111001", 20463 => "11100001", 20465 => "01110011", 20468 => "10001001", 20472 => "00010100", 20474 => "01010011", 20483 => "01110101", 20485 => "11100001", 20487 => "01010111", 20490 => "10111111", 20491 => "10111010", 20496 => "11001101", 20501 => "01100010", 20502 => "10000010", 20503 => "10011110", 20506 => "10111101", 20508 => "10001001", 20509 => "10001001", 20512 => "10110110", 20516 => "11000001", 20517 => "00010000", 20520 => "00111011", 20528 => "01101100", 20529 => "11100000", 20530 => "01011001", 20533 => "00100000", 20534 => "11110000", 20535 => "01010100", 20537 => "00100111", 20540 => "00010000", 20541 => "01000011", 20543 => "11001001", 20544 => "00111000", 20546 => "01000101", 20548 => "10110101", 20549 => "01011000", 20550 => "11100100", 20551 => "11001011", 20553 => "01011001", 20555 => "01011100", 20557 => "01100010", 20558 => "10111100", 20559 => "01101001", 20560 => "01100010", 20562 => "11110011", 20564 => "11110011", 20566 => "01001101", 20567 => "01010101", 20572 => "11000101", 20576 => "11001000", 20577 => "11110000", 20580 => "11101110", 20581 => "10010000", 20583 => "01010111", 20586 => "11111111", 20587 => "11000010", 20588 => "01000011", 20590 => "11010100", 20591 => "00110111", 20594 => "10111011", 20596 => "10011101", 20599 => "10001100", 20601 => "00101100", 20602 => "11001001", 20603 => "10001100", 20604 => "11101101", 20606 => "00100010", 20607 => "10101000", 20608 => "10011000", 20611 => "11110011", 20614 => "11111010", 20616 => "00110111", 20617 => "11100101", 20620 => "11010100", 20623 => "11010001", 20624 => "01100101", 20626 => "00111010", 20630 => "01101110", 20631 => "10001001", 20636 => "10001100", 20637 => "10101110", 20639 => "00110011", 20640 => "11111001", 20641 => "10011000", 20642 => "00111111", 20643 => "00010010", 20644 => "00000101", 20646 => "10111100", 20647 => "10101011", 20648 => "01000101", 20649 => "11000001", 20650 => "11100010", 20651 => "01010110", 20652 => "11100110", 20653 => "11010110", 20654 => "00010011", 20655 => "01010100", 20658 => "11110101", 20659 => "01100100", 20660 => "01010100", 20663 => "11000100", 20664 => "00111010", 20667 => "10100000", 20670 => "10101100", 20672 => "01101011", 20675 => "00011000", 20682 => "11001110", 20688 => "00111001", 20689 => "01010101", 20690 => "11001010", 20691 => "01100011", 20692 => "11010100", 20694 => "00010000", 20697 => "00010100", 20698 => "10110000", 20699 => "01001000", 20702 => "00110011", 20707 => "00000010", 20710 => "01001010", 20711 => "10011101", 20714 => "00100000", 20718 => "01101011", 20720 => "00000101", 20723 => "11100001", 20727 => "00111011", 20731 => "01101010", 20733 => "00101000", 20736 => "00000100", 20737 => "11101111", 20739 => "11111100", 20741 => "10110000", 20742 => "01000100", 20744 => "10001101", 20750 => "11101101", 20751 => "10001010", 20752 => "11010011", 20753 => "00010101", 20758 => "01001101", 20759 => "00001111", 20764 => "11110001", 20767 => "01100010", 20768 => "10001010", 20770 => "00111011", 20771 => "11111000", 20775 => "01010011", 20778 => "11111001", 20780 => "01010001", 20783 => "01110101", 20784 => "10011001", 20789 => "10010100", 20790 => "01011110", 20791 => "01100111", 20792 => "01010010", 20796 => "00000101", 20797 => "10011100", 20798 => "10001100", 20800 => "10001101", 20803 => "00000010", 20804 => "11110001", 20806 => "00010011", 20807 => "00111100", 20810 => "01011110", 20813 => "01100101", 20814 => "10011100", 20816 => "00000111", 20817 => "00110000", 20818 => "01110011", 20825 => "01100101", 20826 => "10010100", 20827 => "10000011", 20828 => "00001111", 20829 => "00000100", 20830 => "00100000", 20831 => "00101010", 20834 => "01000100", 20835 => "01111001", 20838 => "10001101", 20840 => "11100110", 20841 => "01100100", 20843 => "00111110", 20845 => "10101010", 20848 => "01001001", 20850 => "11011011", 20853 => "01110101", 20854 => "11101001", 20855 => "01111000", 20857 => "00001111", 20864 => "10010011", 20867 => "01111101", 20868 => "11001001", 20869 => "10010010", 20871 => "01010010", 20875 => "00100001", 20877 => "11001110", 20879 => "01000000", 20880 => "00001100", 20881 => "11101010", 20882 => "11011010", 20884 => "10100011", 20889 => "00101010", 20890 => "00100001", 20894 => "11110000", 20897 => "11010111", 20900 => "00101111", 20901 => "00000110", 20903 => "01001011", 20904 => "01010101", 20905 => "01011100", 20906 => "11100111", 20907 => "00110100", 20908 => "00100001", 20909 => "00100000", 20910 => "11001010", 20911 => "01000001", 20914 => "00101101", 20917 => "11011110", 20918 => "00001000", 20921 => "00011111", 20922 => "10100110", 20925 => "10001111", 20927 => "01110100", 20932 => "00111111", 20933 => "00001010", 20935 => "11110001", 20936 => "01011000", 20938 => "01111100", 20940 => "00010000", 20941 => "00111111", 20942 => "11110011", 20943 => "01111101", 20946 => "11010100", 20947 => "00110100", 20949 => "11111110", 20952 => "11011100", 20955 => "10000000", 20957 => "01111011", 20958 => "01010100", 20960 => "11001111", 20964 => "00010011", 20967 => "11110101", 20968 => "01010101", 20969 => "01001100", 20971 => "00011010", 20972 => "01100101", 20973 => "11011011", 20977 => "10110010", 20978 => "11010001", 20979 => "01110111", 20980 => "10110000", 20982 => "11111111", 20984 => "10101110", 20987 => "10100110", 20989 => "11101011", 20991 => "10000110", 20993 => "01101100", 20995 => "01011111", 21000 => "11100101", 21001 => "01100100", 21003 => "11101101", 21004 => "11100100", 21006 => "00001011", 21008 => "00010100", 21012 => "10011001", 21013 => "10001100", 21017 => "00010110", 21019 => "01100110", 21030 => "10010000", 21033 => "10100001", 21038 => "11110001", 21039 => "11101100", 21040 => "10011010", 21042 => "11110110", 21043 => "11001010", 21044 => "00001100", 21045 => "01111000", 21047 => "10011111", 21049 => "11111111", 21051 => "11100001", 21053 => "01000011", 21055 => "11010101", 21058 => "00101100", 21061 => "10011110", 21064 => "01001000", 21065 => "00001110", 21066 => "11000011", 21067 => "00011100", 21068 => "00110001", 21070 => "00100000", 21071 => "11100011", 21072 => "01010000", 21073 => "11010101", 21074 => "10111000", 21077 => "11011001", 21078 => "11001000", 21084 => "10000011", 21089 => "11100110", 21090 => "01001111", 21091 => "00010101", 21095 => "01111011", 21100 => "00001010", 21103 => "01001011", 21106 => "01000001", 21110 => "01100011", 21111 => "10010010", 21112 => "11110001", 21113 => "00110011", 21114 => "00100100", 21116 => "11010100", 21117 => "10110001", 21118 => "10000001", 21120 => "11001100", 21126 => "10100101", 21128 => "10011110", 21130 => "10110111", 21131 => "10010000", 21136 => "11011101", 21138 => "01011101", 21141 => "10011001", 21142 => "11011011", 21144 => "01101010", 21147 => "10110111", 21148 => "10011011", 21150 => "00000101", 21152 => "10001110", 21154 => "00100100", 21155 => "00000011", 21158 => "01000100", 21159 => "11000111", 21163 => "11100111", 21168 => "01011101", 21169 => "11111100", 21170 => "11000100", 21173 => "01000110", 21174 => "10111010", 21176 => "10101000", 21177 => "01011111", 21180 => "00101110", 21181 => "01010011", 21182 => "01010001", 21183 => "01011000", 21185 => "10011001", 21189 => "10001011", 21190 => "11100111", 21191 => "00010100", 21192 => "01101000", 21194 => "00100110", 21195 => "10000101", 21196 => "00101101", 21197 => "11100011", 21198 => "00000110", 21200 => "01011111", 21202 => "11111110", 21203 => "10000011", 21204 => "11110101", 21205 => "10011011", 21206 => "10111001", 21208 => "10101000", 21209 => "11111100", 21211 => "11001000", 21215 => "10111001", 21216 => "00000111", 21217 => "10101011", 21218 => "11101110", 21219 => "11100010", 21220 => "11111000", 21221 => "01000111", 21223 => "00111111", 21224 => "01111111", 21227 => "00110101", 21228 => "10000010", 21230 => "00101001", 21232 => "11111000", 21233 => "10111001", 21234 => "00010010", 21239 => "01011101", 21241 => "10100110", 21244 => "00111101", 21245 => "11100001", 21248 => "01010011", 21250 => "10111001", 21253 => "01111111", 21254 => "11000101", 21259 => "01001000", 21260 => "11010001", 21263 => "11001101", 21266 => "00011011", 21269 => "11000011", 21271 => "00110110", 21272 => "10001111", 21274 => "01101011", 21276 => "01011001", 21278 => "00000100", 21279 => "01001000", 21283 => "01111011", 21287 => "10111111", 21289 => "10001011", 21293 => "00101100", 21295 => "00010111", 21296 => "11101011", 21297 => "01011000", 21299 => "01100110", 21304 => "01100001", 21305 => "00100100", 21306 => "10001111", 21308 => "01111101", 21309 => "01101001", 21311 => "11100111", 21315 => "00110011", 21316 => "00100110", 21317 => "11111101", 21318 => "01111111", 21319 => "01111111", 21323 => "10101111", 21328 => "10110111", 21331 => "10001010", 21332 => "00100000", 21333 => "10001001", 21336 => "01000100", 21340 => "10000110", 21344 => "11100110", 21345 => "00010101", 21346 => "01011100", 21347 => "01100111", 21348 => "01100000", 21354 => "00111101", 21355 => "01110100", 21358 => "00110010", 21361 => "01001111", 21363 => "01011001", 21368 => "00110110", 21369 => "10001110", 21370 => "11100101", 21373 => "11001011", 21376 => "10100101", 21377 => "01110000", 21379 => "00011111", 21380 => "01010111", 21382 => "01110100", 21383 => "11001101", 21388 => "01011110", 21390 => "11010010", 21394 => "00110101", 21398 => "11010101", 21399 => "10100000", 21400 => "01011100", 21401 => "10111100", 21404 => "00100100", 21406 => "00111110", 21409 => "10000110", 21411 => "01010001", 21414 => "00010001", 21415 => "00001101", 21416 => "00000111", 21421 => "01101100", 21423 => "11011100", 21424 => "01011100", 21425 => "11001011", 21426 => "00100010", 21428 => "10001110", 21431 => "01001101", 21435 => "01001111", 21436 => "01110011", 21438 => "01001000", 21444 => "01011000", 21446 => "11010101", 21448 => "11110100", 21449 => "11110000", 21451 => "11100101", 21457 => "01111000", 21461 => "01110001", 21462 => "00111001", 21466 => "10110111", 21467 => "10100010", 21469 => "01001110", 21470 => "01110100", 21472 => "11010001", 21474 => "11010101", 21476 => "00100110", 21477 => "10101110", 21479 => "00010110", 21480 => "11010000", 21482 => "11101011", 21484 => "00101110", 21488 => "11111010", 21489 => "00110101", 21490 => "11110000", 21492 => "11001100", 21493 => "11010111", 21494 => "10101100", 21499 => "10101110", 21501 => "11101111", 21502 => "00111011", 21503 => "10111011", 21504 => "00000110", 21505 => "10011000", 21506 => "00011011", 21507 => "01110100", 21508 => "11010101", 21512 => "01010100", 21514 => "00101101", 21517 => "01111110", 21520 => "01111011", 21526 => "11000010", 21536 => "11101111", 21538 => "01110000", 21539 => "11111100", 21541 => "10101001", 21542 => "01011001", 21545 => "11101100", 21547 => "11010000", 21550 => "11010011", 21553 => "01100100", 21557 => "00111111", 21558 => "00110001", 21560 => "01100001", 21561 => "11100011", 21562 => "01110000", 21572 => "11110000", 21574 => "10100000", 21576 => "10000100", 21577 => "10011111", 21578 => "00000100", 21579 => "11011011", 21585 => "10010111", 21587 => "10100011", 21589 => "11100000", 21590 => "10101010", 21591 => "01101001", 21592 => "10011101", 21593 => "00101010", 21594 => "00111111", 21595 => "10100000", 21596 => "10100010", 21597 => "01110011", 21598 => "01110110", 21599 => "10111100", 21607 => "00100100", 21609 => "10101110", 21610 => "10110110", 21612 => "11001010", 21613 => "10001110", 21615 => "01100010", 21616 => "11001100", 21617 => "00010100", 21618 => "00101101", 21621 => "11000101", 21624 => "01001101", 21625 => "01101111", 21629 => "00111101", 21631 => "11011110", 21632 => "00011001", 21633 => "01000101", 21636 => "01101000", 21640 => "11111011", 21641 => "11101000", 21642 => "01111001", 21644 => "01111010", 21645 => "10111010", 21647 => "01110010", 21648 => "11110110", 21650 => "11110101", 21651 => "10011001", 21653 => "00110111", 21654 => "00001011", 21658 => "01100100", 21659 => "11111000", 21664 => "10010001", 21667 => "01111110", 21669 => "10110111", 21670 => "10110011", 21672 => "11100001", 21675 => "01111001", 21677 => "00010110", 21682 => "01100101", 21685 => "01110111", 21687 => "00010100", 21689 => "01000010", 21695 => "01011001", 21701 => "11010011", 21703 => "00010001", 21704 => "00000010", 21705 => "00100101", 21706 => "10101101", 21707 => "01100110", 21709 => "00110110", 21711 => "10011100", 21712 => "01000100", 21713 => "10011001", 21717 => "11110000", 21720 => "01110101", 21721 => "10000101", 21723 => "01001000", 21725 => "10100010", 21728 => "00100001", 21730 => "01100001", 21731 => "00101011", 21734 => "01011011", 21736 => "11011000", 21737 => "00001101", 21738 => "00111000", 21739 => "00111101", 21741 => "00011111", 21744 => "00101000", 21746 => "10001100", 21747 => "00101110", 21749 => "01011011", 21753 => "01011000", 21755 => "01101001", 21756 => "01000011", 21757 => "00101100", 21759 => "01001100", 21760 => "00110010", 21762 => "00000010", 21764 => "10100100", 21765 => "10101001", 21768 => "01111001", 21773 => "10110000", 21774 => "10000010", 21777 => "01010111", 21779 => "10100000", 21783 => "00001101", 21784 => "01000110", 21785 => "01100100", 21788 => "11100110", 21790 => "00001100", 21792 => "00111001", 21793 => "11111010", 21797 => "10110110", 21799 => "11110111", 21802 => "00100100", 21803 => "01111101", 21804 => "00111011", 21808 => "01101100", 21811 => "10111111", 21814 => "01000101", 21815 => "11011100", 21818 => "00011011", 21819 => "01101000", 21820 => "00100001", 21826 => "11101110", 21827 => "01100110", 21830 => "00100011", 21832 => "11001100", 21833 => "10110001", 21834 => "01111000", 21836 => "01110110", 21838 => "01001000", 21839 => "11010011", 21841 => "01010010", 21844 => "11100101", 21847 => "11001111", 21850 => "00010101", 21853 => "01000011", 21854 => "10100101", 21855 => "10101111", 21861 => "00101011", 21865 => "10110100", 21866 => "01011010", 21868 => "00111110", 21872 => "01101011", 21873 => "11001110", 21874 => "10100100", 21875 => "10010001", 21878 => "11111100", 21885 => "11001110", 21887 => "10110110", 21888 => "11110100", 21889 => "10001010", 21890 => "10111011", 21891 => "01011111", 21892 => "01100001", 21893 => "11010111", 21897 => "10101010", 21899 => "10101100", 21901 => "00110100", 21903 => "01101011", 21905 => "11010001", 21908 => "00100001", 21909 => "00011100", 21910 => "00100100", 21913 => "01001001", 21920 => "11100110", 21922 => "11000011", 21925 => "11100000", 21927 => "11101001", 21930 => "01100001", 21932 => "10000011", 21936 => "01001100", 21937 => "11110000", 21941 => "10100101", 21943 => "00011000", 21946 => "11100010", 21950 => "00001001", 21952 => "00110001", 21953 => "10111001", 21954 => "00100011", 21957 => "11011100", 21958 => "00101000", 21959 => "00111011", 21961 => "11000110", 21964 => "00101100", 21966 => "11101100", 21967 => "10000100", 21968 => "01110000", 21970 => "01100000", 21972 => "11010110", 21978 => "00111010", 21979 => "11000100", 21980 => "01100110", 21981 => "10100000", 21985 => "11000111", 21986 => "01111010", 21987 => "01100111", 21989 => "00110110", 21995 => "00110110", 21996 => "10010100", 21999 => "10111111", 22002 => "11011011", 22006 => "00111001", 22007 => "01001010", 22012 => "00001010", 22013 => "01010111", 22014 => "10000011", 22015 => "00010111", 22020 => "01101101", 22021 => "00000010", 22022 => "00010110", 22025 => "00001110", 22026 => "01011000", 22028 => "10000010", 22031 => "00011101", 22032 => "10000001", 22033 => "00101010", 22034 => "10101101", 22035 => "00101010", 22036 => "10001100", 22037 => "01110000", 22038 => "01001110", 22040 => "11010000", 22041 => "10101001", 22043 => "10010001", 22044 => "11010111", 22046 => "10100100", 22047 => "01010001", 22049 => "01000001", 22050 => "11011011", 22052 => "11110101", 22053 => "00100101", 22054 => "01011110", 22057 => "01011101", 22058 => "11010011", 22063 => "01010011", 22066 => "10010011", 22067 => "11000011", 22068 => "01011101", 22074 => "00000011", 22075 => "10011000", 22080 => "11000000", 22081 => "00101010", 22084 => "11110001", 22085 => "11110010", 22086 => "00100011", 22087 => "10010101", 22091 => "00001011", 22097 => "10101010", 22098 => "11011111", 22100 => "00011000", 22101 => "11011111", 22102 => "10110010", 22104 => "10101111", 22105 => "01111001", 22106 => "01000000", 22107 => "11011101", 22108 => "01111100", 22112 => "00000010", 22114 => "00001101", 22117 => "10111111", 22119 => "10001110", 22120 => "01100100", 22121 => "00001011", 22123 => "01110100", 22126 => "00001100", 22131 => "01101100", 22132 => "01011001", 22137 => "01000110", 22142 => "11111000", 22144 => "01010010", 22147 => "01010011", 22148 => "01001111", 22150 => "11100010", 22152 => "11101000", 22154 => "00010001", 22159 => "00111100", 22161 => "00001100", 22163 => "00001110", 22164 => "10011101", 22166 => "00100101", 22167 => "11010100", 22168 => "11100010", 22171 => "11110001", 22172 => "01100100", 22178 => "10101000", 22179 => "10010100", 22182 => "11111100", 22184 => "10111011", 22189 => "01001000", 22190 => "10111010", 22193 => "11011010", 22195 => "00110010", 22196 => "10010110", 22197 => "10000100", 22199 => "11110110", 22201 => "01101001", 22203 => "10100101", 22207 => "10110010", 22208 => "00010101", 22212 => "11110100", 22213 => "00000010", 22214 => "10110010", 22218 => "10000111", 22219 => "00111000", 22222 => "00100110", 22223 => "00111010", 22231 => "01100110", 22232 => "01010010", 22242 => "11001100", 22244 => "01100000", 22249 => "10000100", 22251 => "11000001", 22252 => "11101011", 22253 => "10000101", 22254 => "01101111", 22255 => "01110000", 22257 => "11011110", 22258 => "10101100", 22259 => "10000000", 22260 => "00000101", 22264 => "10000101", 22265 => "01011110", 22268 => "10010011", 22270 => "00001111", 22273 => "11110000", 22275 => "01010010", 22280 => "01010111", 22281 => "00011111", 22282 => "10110011", 22284 => "01111010", 22292 => "01001010", 22293 => "11101100", 22297 => "01010100", 22299 => "00111011", 22301 => "10101001", 22306 => "01111000", 22310 => "00111001", 22311 => "10100101", 22315 => "00100001", 22318 => "00111111", 22320 => "10100101", 22324 => "11000010", 22327 => "10110000", 22332 => "11011001", 22333 => "00010000", 22334 => "00100011", 22335 => "10111010", 22336 => "11111010", 22337 => "11110010", 22339 => "11101011", 22342 => "10010001", 22346 => "00110110", 22347 => "11010000", 22348 => "11011110", 22351 => "01100000", 22354 => "11110001", 22357 => "11011011", 22358 => "11111111", 22359 => "10011010", 22361 => "11000011", 22365 => "01101111", 22366 => "01101111", 22368 => "00000110", 22369 => "00011101", 22375 => "10001001", 22376 => "11011111", 22377 => "01111011", 22378 => "10110000", 22380 => "01001111", 22382 => "01001101", 22383 => "01011101", 22386 => "01100101", 22388 => "11101001", 22389 => "00101001", 22390 => "01010011", 22394 => "01000001", 22408 => "10101111", 22411 => "01110111", 22412 => "10001100", 22414 => "01101001", 22415 => "10111110", 22417 => "00111000", 22418 => "10010011", 22419 => "00010111", 22420 => "10101100", 22422 => "01001000", 22424 => "11111000", 22425 => "10111101", 22426 => "10100010", 22427 => "10011110", 22430 => "10101000", 22431 => "11100011", 22432 => "00101101", 22433 => "11111011", 22434 => "10001000", 22435 => "00111111", 22436 => "10000011", 22440 => "00111101", 22444 => "01110111", 22446 => "00111001", 22447 => "00101011", 22450 => "10110101", 22451 => "10001101", 22452 => "01010110", 22453 => "01100010", 22454 => "10111011", 22456 => "00011110", 22458 => "00011101", 22459 => "10001101", 22460 => "11110011", 22461 => "01110001", 22465 => "00110110", 22466 => "00111110", 22467 => "00101010", 22470 => "01100010", 22472 => "00010001", 22474 => "11001001", 22476 => "01110011", 22477 => "10100011", 22478 => "10000111", 22485 => "01110011", 22487 => "10010001", 22489 => "01010010", 22492 => "11010000", 22494 => "00000011", 22496 => "01001110", 22500 => "10001110", 22501 => "01001011", 22502 => "11000001", 22504 => "01000100", 22506 => "01011101", 22507 => "00001111", 22508 => "00010100", 22510 => "10000101", 22512 => "01011100", 22513 => "00001101", 22521 => "00100110", 22524 => "10011101", 22530 => "00011011", 22531 => "00110111", 22533 => "10111101", 22535 => "10101110", 22538 => "10100110", 22539 => "11111110", 22542 => "11110100", 22545 => "11111000", 22551 => "11111111", 22554 => "01100001", 22556 => "11000100", 22558 => "11111110", 22560 => "00001001", 22561 => "01110001", 22564 => "00100001", 22565 => "10101011", 22566 => "01010100", 22569 => "00111110", 22574 => "00100100", 22579 => "01100001", 22582 => "10001001", 22583 => "01010111", 22587 => "10101100", 22590 => "00100100", 22591 => "01010101", 22592 => "01100011", 22595 => "00100000", 22600 => "11100000", 22606 => "10101011", 22608 => "11001001", 22611 => "10101111", 22613 => "11100011", 22617 => "01111100", 22619 => "01011100", 22621 => "01101111", 22622 => "11111110", 22624 => "01000111", 22627 => "11100011", 22628 => "10111111", 22631 => "00011000", 22633 => "01111100", 22635 => "01111010", 22636 => "00011111", 22637 => "11100110", 22638 => "10010011", 22640 => "01100011", 22644 => "00011101", 22645 => "11000110", 22649 => "00111101", 22650 => "10011111", 22653 => "11101100", 22654 => "00110010", 22655 => "00110001", 22656 => "00100000", 22660 => "00101000", 22666 => "00001111", 22668 => "00000111", 22671 => "10111110", 22673 => "01011000", 22676 => "11011101", 22679 => "11100110", 22682 => "10001100", 22684 => "10011011", 22685 => "11110110", 22690 => "01000010", 22695 => "01101101", 22697 => "11011111", 22698 => "01101011", 22700 => "00111001", 22701 => "11001001", 22703 => "00001110", 22704 => "00100101", 22705 => "11110111", 22708 => "00110110", 22710 => "10001111", 22711 => "01101000", 22715 => "10101111", 22716 => "10111011", 22720 => "00000101", 22721 => "10111001", 22724 => "00001100", 22725 => "01101110", 22727 => "11110101", 22729 => "10101110", 22731 => "11010011", 22732 => "01001001", 22739 => "00010011", 22740 => "10000111", 22741 => "11010111", 22743 => "10010001", 22744 => "01110110", 22748 => "00001011", 22751 => "01100010", 22753 => "11100000", 22758 => "01100100", 22760 => "00111000", 22761 => "11100010", 22764 => "11110100", 22765 => "00000100", 22767 => "01000110", 22769 => "01110010", 22771 => "01100110", 22772 => "10001001", 22773 => "01001010", 22774 => "11110000", 22775 => "01010100", 22777 => "01010110", 22778 => "11010100", 22779 => "01000110", 22780 => "11010000", 22783 => "00011001", 22785 => "11110001", 22786 => "00111010", 22787 => "11101011", 22788 => "01111011", 22789 => "11000010", 22790 => "01001101", 22791 => "01010010", 22795 => "10111011", 22798 => "01101010", 22800 => "10000110", 22801 => "00011100", 22804 => "10100010", 22805 => "11101110", 22807 => "01110010", 22808 => "00110110", 22812 => "11110010", 22815 => "11000001", 22819 => "00001111", 22821 => "01100110", 22822 => "01111011", 22825 => "00010010", 22829 => "10000001", 22830 => "00111011", 22831 => "00010001", 22832 => "10111000", 22835 => "00110101", 22836 => "11100010", 22838 => "00100111", 22841 => "00000110", 22842 => "00110000", 22844 => "01011011", 22846 => "11001001", 22848 => "00001100", 22853 => "10110111", 22858 => "00010000", 22859 => "00110100", 22860 => "01101101", 22861 => "11011000", 22864 => "10101011", 22865 => "11111100", 22866 => "10011111", 22867 => "00101110", 22868 => "10111111", 22869 => "00100001", 22870 => "10010101", 22872 => "00110101", 22874 => "00110111", 22876 => "01100101", 22879 => "11111101", 22880 => "00101110", 22881 => "00110000", 22882 => "11111001", 22883 => "10111010", 22886 => "01010100", 22887 => "10011011", 22888 => "11100110", 22889 => "01001110", 22893 => "01010101", 22894 => "10010000", 22899 => "01101111", 22904 => "10100110", 22905 => "01110111", 22906 => "10000010", 22907 => "10100111", 22908 => "00000011", 22913 => "00001111", 22918 => "10011000", 22923 => "00000001", 22928 => "10010001", 22929 => "00011011", 22932 => "11110101", 22937 => "01000001", 22939 => "10110011", 22943 => "11001011", 22945 => "00101001", 22947 => "00100110", 22949 => "00000010", 22952 => "01010101", 22953 => "01011010", 22956 => "10100010", 22958 => "00110001", 22959 => "11100011", 22960 => "10011110", 22961 => "10000011", 22962 => "10100100", 22963 => "01111010", 22964 => "11001100", 22967 => "00001001", 22971 => "11110101", 22974 => "00011110", 22975 => "01001110", 22977 => "10101010", 22979 => "00010010", 22980 => "10001000", 22983 => "01000010", 22984 => "10001110", 22985 => "11101001", 22988 => "01101111", 22989 => "11011100", 22993 => "11011001", 22994 => "01001000", 22995 => "10010110", 22996 => "01000100", 23001 => "00001000", 23002 => "01100100", 23004 => "10001010", 23005 => "10001000", 23006 => "11100101", 23010 => "00111001", 23013 => "10011000", 23014 => "01011010", 23017 => "11100001", 23018 => "00110100", 23019 => "01101101", 23020 => "01011100", 23021 => "11101100", 23023 => "10101101", 23024 => "01100110", 23025 => "00100001", 23026 => "10011100", 23027 => "00011001", 23029 => "10110110", 23030 => "10110101", 23032 => "01001110", 23034 => "10010100", 23035 => "11000111", 23037 => "00001111", 23038 => "10001011", 23039 => "11000110", 23040 => "10010011", 23042 => "10001110", 23043 => "01111111", 23045 => "01100110", 23050 => "11010111", 23053 => "00111011", 23057 => "11001001", 23058 => "11001101", 23060 => "10101111", 23061 => "11100011", 23062 => "00111100", 23064 => "01111001", 23065 => "00001001", 23067 => "10111101", 23068 => "00000100", 23072 => "00010111", 23074 => "10101000", 23076 => "11011110", 23078 => "11010111", 23079 => "11011110", 23081 => "01110010", 23084 => "10101001", 23087 => "10010101", 23088 => "10001101", 23089 => "01001001", 23090 => "10001111", 23091 => "01111101", 23092 => "11011110", 23094 => "10110110", 23095 => "10101001", 23096 => "10111011", 23098 => "01011110", 23099 => "01110101", 23100 => "10001001", 23103 => "10100110", 23108 => "10011101", 23109 => "11100011", 23110 => "10001111", 23111 => "11100001", 23114 => "10000010", 23118 => "11010100", 23119 => "10100111", 23120 => "00110110", 23121 => "10110101", 23122 => "00110011", 23123 => "11100001", 23125 => "10001110", 23126 => "11011001", 23127 => "11111001", 23128 => "11111111", 23132 => "10000010", 23134 => "10000010", 23137 => "11101010", 23140 => "01101100", 23141 => "00111011", 23142 => "00011101", 23147 => "01110111", 23149 => "00000111", 23150 => "11100010", 23153 => "10000001", 23155 => "10101011", 23157 => "00011011", 23159 => "11001010", 23160 => "01100010", 23163 => "01100000", 23164 => "01011101", 23167 => "11110101", 23168 => "11001101", 23171 => "01101011", 23172 => "11111110", 23174 => "01001110", 23175 => "01000001", 23179 => "11110101", 23180 => "01100011", 23183 => "10001000", 23184 => "10100011", 23185 => "11101101", 23186 => "11110001", 23189 => "01000000", 23191 => "01100000", 23192 => "10101111", 23196 => "10001110", 23199 => "10100000", 23200 => "00110101", 23204 => "00110100", 23206 => "11010101", 23207 => "01010010", 23209 => "11001000", 23210 => "11101100", 23211 => "10110101", 23212 => "11001001", 23213 => "10001100", 23219 => "10101111", 23220 => "01101111", 23221 => "01100001", 23224 => "01000101", 23225 => "10010010", 23227 => "10101110", 23228 => "01000010", 23231 => "01110101", 23232 => "01110010", 23246 => "10010100", 23249 => "10001110", 23250 => "01111011", 23251 => "00000110", 23253 => "01101010", 23254 => "11011111", 23259 => "10100010", 23261 => "00000111", 23263 => "00111001", 23264 => "11101010", 23265 => "01011101", 23267 => "01001110", 23273 => "11001101", 23274 => "01011101", 23276 => "11101001", 23277 => "00011111", 23280 => "00001111", 23282 => "11101000", 23283 => "10010110", 23285 => "10111111", 23286 => "11000000", 23290 => "00101100", 23296 => "11101001", 23298 => "01111000", 23299 => "00001110", 23300 => "11011001", 23302 => "11101100", 23303 => "01011111", 23304 => "00000110", 23306 => "11101101", 23307 => "11011101", 23310 => "11101100", 23318 => "01011001", 23319 => "01000101", 23320 => "10011001", 23322 => "00100000", 23323 => "11001110", 23326 => "01100101", 23327 => "11110001", 23328 => "10010010", 23335 => "11001010", 23342 => "00110001", 23345 => "00101001", 23346 => "10100111", 23350 => "01101010", 23355 => "01011000", 23358 => "10001100", 23360 => "00110110", 23363 => "11101101", 23364 => "10011110", 23365 => "10100011", 23367 => "01000011", 23368 => "11111000", 23369 => "10101010", 23374 => "00110100", 23375 => "01111110", 23377 => "10001111", 23380 => "00111110", 23383 => "10110110", 23385 => "10111011", 23386 => "00111001", 23387 => "01101110", 23389 => "00001110", 23390 => "11110000", 23391 => "01101011", 23393 => "10110111", 23394 => "01000111", 23395 => "00000001", 23396 => "01111100", 23397 => "11000110", 23398 => "00110101", 23403 => "01111110", 23406 => "00000011", 23407 => "00100101", 23409 => "10011101", 23410 => "01000010", 23411 => "10100101", 23412 => "00101110", 23413 => "01111000", 23414 => "11111111", 23415 => "01000101", 23416 => "11101111", 23417 => "10100100", 23418 => "11110100", 23419 => "01000010", 23422 => "00101000", 23424 => "10101011", 23427 => "11010110", 23428 => "11100000", 23429 => "00001101", 23430 => "10100110", 23432 => "10011010", 23433 => "11111100", 23436 => "11001000", 23440 => "00111000", 23441 => "00010100", 23442 => "00110010", 23443 => "11001001", 23444 => "00110101", 23447 => "11000000", 23449 => "11010101", 23450 => "10100101", 23451 => "11111101", 23452 => "10011111", 23460 => "00010001", 23463 => "00100000", 23464 => "10101010", 23465 => "10010110", 23470 => "10000000", 23471 => "01111111", 23473 => "00001100", 23474 => "01001110", 23477 => "01001101", 23478 => "10111001", 23481 => "10001000", 23482 => "01010001", 23483 => "10111011", 23486 => "00010111", 23489 => "10010010", 23493 => "00011000", 23495 => "11010101", 23496 => "00111010", 23497 => "11110011", 23502 => "00010001", 23503 => "10010000", 23504 => "11010001", 23505 => "00100110", 23507 => "10010100", 23511 => "00101001", 23512 => "11010011", 23514 => "01000001", 23515 => "01001001", 23518 => "01001011", 23521 => "00000001", 23522 => "10010101", 23523 => "11101111", 23524 => "01111010", 23526 => "00011101", 23530 => "10101100", 23532 => "01000101", 23535 => "01010001", 23539 => "00010001", 23543 => "10011010", 23544 => "01000011", 23547 => "11111100", 23549 => "00000011", 23555 => "00101000", 23557 => "00101010", 23558 => "01101001", 23559 => "10111000", 23560 => "10000011", 23567 => "11000010", 23569 => "11111011", 23570 => "11000011", 23572 => "01000110", 23573 => "00001001", 23574 => "01011011", 23575 => "00100010", 23576 => "11001100", 23577 => "01111010", 23578 => "10011010", 23584 => "00001011", 23585 => "01000000", 23586 => "00100100", 23587 => "00001101", 23589 => "00110111", 23590 => "10011100", 23591 => "00101000", 23595 => "10001100", 23596 => "11001001", 23597 => "10110110", 23598 => "11001101", 23599 => "11100101", 23602 => "01011000", 23603 => "01000001", 23604 => "10100111", 23605 => "00001011", 23606 => "00100101", 23608 => "00001100", 23610 => "01101101", 23611 => "10101010", 23612 => "10000110", 23615 => "00000101", 23616 => "11111010", 23620 => "11010100", 23621 => "01000100", 23622 => "10010010", 23623 => "11010111", 23625 => "00001101", 23627 => "11111011", 23628 => "10111111", 23629 => "10100000", 23631 => "11000010", 23632 => "00110010", 23637 => "00101011", 23638 => "10100111", 23639 => "01010101", 23641 => "01000001", 23642 => "00010010", 23643 => "01010010", 23644 => "11110010", 23650 => "01111110", 23651 => "11011100", 23652 => "11110110", 23653 => "01111000", 23658 => "10111111", 23660 => "11101001", 23662 => "00110100", 23663 => "11001000", 23671 => "11100001", 23673 => "11110100", 23675 => "11011101", 23676 => "11100100", 23679 => "00000100", 23680 => "11110100", 23682 => "11111111", 23685 => "10111000", 23686 => "00111000", 23689 => "11000010", 23690 => "00110111", 23691 => "00010100", 23693 => "00100110", 23701 => "01010010", 23707 => "11101110", 23710 => "11011010", 23712 => "01011010", 23713 => "11111101", 23715 => "11000101", 23717 => "10010000", 23719 => "00010010", 23723 => "01001101", 23726 => "10111000", 23728 => "11001110", 23729 => "00011011", 23732 => "00111101", 23733 => "00111110", 23734 => "10001010", 23735 => "10101100", 23736 => "10010010", 23738 => "11001101", 23739 => "10011100", 23740 => "11001001", 23742 => "01001011", 23743 => "11000100", 23745 => "00101000", 23746 => "01100000", 23747 => "10011010", 23748 => "11101110", 23751 => "11011001", 23752 => "01101101", 23755 => "10001111", 23757 => "10100111", 23762 => "00000100", 23763 => "01110001", 23768 => "00110111", 23769 => "01010001", 23773 => "10001011", 23774 => "10111001", 23775 => "00100101", 23780 => "10011011", 23784 => "11000111", 23785 => "11000010", 23789 => "11101100", 23790 => "01010110", 23791 => "01011011", 23792 => "10111111", 23795 => "11110010", 23797 => "10110010", 23798 => "11001000", 23802 => "01110101", 23803 => "01001001", 23804 => "10000111", 23805 => "10011101", 23809 => "00011011", 23812 => "01011010", 23813 => "10011101", 23814 => "10100001", 23815 => "01100100", 23819 => "00100010", 23820 => "00011011", 23821 => "00110100", 23823 => "01010001", 23825 => "00000011", 23829 => "11110001", 23832 => "01001101", 23836 => "10001101", 23838 => "00001110", 23841 => "01011001", 23842 => "10100001", 23843 => "01101011", 23844 => "00110111", 23846 => "11000001", 23847 => "11111011", 23848 => "01010110", 23850 => "01011010", 23851 => "10000011", 23854 => "11001000", 23855 => "00000101", 23857 => "01011001", 23860 => "10001110", 23864 => "10101111", 23865 => "10101010", 23867 => "11001111", 23869 => "00110110", 23870 => "11110111", 23872 => "10010110", 23875 => "00110001", 23877 => "01000001", 23884 => "00110001", 23888 => "01111010", 23889 => "00011100", 23890 => "10000101", 23892 => "01101101", 23894 => "01111001", 23901 => "01000111", 23904 => "10100100", 23908 => "00001101", 23913 => "00101100", 23914 => "11010001", 23915 => "10010010", 23916 => "10101111", 23917 => "11111000", 23918 => "11111111", 23920 => "11010100", 23925 => "11000111", 23928 => "00010000", 23929 => "01111101", 23938 => "01100110", 23939 => "11100101", 23940 => "10110111", 23942 => "01111101", 23945 => "00101011", 23948 => "01010001", 23952 => "01101110", 23953 => "01101001", 23955 => "10101110", 23956 => "10110000", 23959 => "01111011", 23962 => "01011111", 23963 => "11010110", 23964 => "01111110", 23965 => "10101100", 23967 => "10011101", 23971 => "00011010", 23972 => "00100001", 23973 => "00111001", 23974 => "11000000", 23975 => "00100110", 23976 => "10001101", 23981 => "01011101", 23983 => "01010101", 23986 => "01110011", 23987 => "00111100", 23993 => "11010010", 23996 => "01101101", 23997 => "00110011", 23998 => "00011000", 23999 => "11110100", 24004 => "00000011", 24010 => "10011001", 24012 => "01001011", 24017 => "00010111", 24019 => "11100101", 24020 => "00000011", 24021 => "00010100", 24025 => "01111001", 24028 => "01001111", 24029 => "00011110", 24031 => "00001001", 24040 => "01010010", 24042 => "01000111", 24043 => "01111011", 24044 => "11000100", 24045 => "10010001", 24051 => "00101010", 24052 => "11101010", 24053 => "11101100", 24054 => "10101101", 24056 => "11011010", 24057 => "10110000", 24058 => "11100000", 24059 => "01010100", 24061 => "01110010", 24063 => "00110101", 24066 => "10011011", 24070 => "01001101", 24074 => "00101001", 24075 => "00000010", 24077 => "11110101", 24078 => "00011100", 24079 => "00110000", 24080 => "00000010", 24081 => "11010011", 24084 => "11010111", 24085 => "01101110", 24089 => "01001100", 24090 => "10010001", 24095 => "11011010", 24096 => "10010011", 24098 => "00100011", 24099 => "01001110", 24104 => "00000111", 24105 => "00010000", 24106 => "11100011", 24107 => "00000010", 24108 => "00101001", 24109 => "10100110", 24110 => "00001111", 24112 => "11000110", 24114 => "00101001", 24115 => "00010010", 24123 => "10000001", 24126 => "10011100", 24129 => "00101001", 24130 => "11011101", 24131 => "11010000", 24132 => "01111110", 24133 => "00101110", 24135 => "00100111", 24137 => "00011010", 24138 => "00110111", 24140 => "01010111", 24141 => "00100010", 24143 => "00000110", 24144 => "11110010", 24146 => "11010110", 24147 => "11010101", 24152 => "10001010", 24154 => "11111000", 24155 => "01110011", 24156 => "11100011", 24158 => "00011101", 24159 => "00010100", 24160 => "00011001", 24162 => "01000111", 24165 => "01011001", 24169 => "01100001", 24170 => "11010010", 24171 => "01010100", 24172 => "00100111", 24176 => "10010000", 24180 => "10000011", 24186 => "11011001", 24187 => "10111111", 24188 => "00100101", 24190 => "11011110", 24192 => "11000001", 24193 => "00110110", 24196 => "00110111", 24198 => "11110101", 24201 => "00111110", 24203 => "11010001", 24205 => "01110001", 24211 => "11001010", 24212 => "10101001", 24214 => "00001111", 24220 => "11101100", 24222 => "00010101", 24225 => "11111111", 24226 => "00101011", 24228 => "11001000", 24229 => "11101001", 24234 => "10011000", 24235 => "00100111", 24236 => "00110000", 24238 => "11000000", 24240 => "11001010", 24241 => "01000101", 24245 => "11111001", 24247 => "00101110", 24248 => "10111010", 24249 => "10010100", 24251 => "00000100", 24260 => "11001001", 24262 => "10100011", 24267 => "01101001", 24270 => "00001101", 24271 => "10010000", 24272 => "01000001", 24273 => "11111010", 24276 => "10011101", 24277 => "11011100", 24280 => "01001101", 24281 => "10000111", 24282 => "11101000", 24285 => "11110001", 24286 => "00100010", 24287 => "11011001", 24288 => "10111111", 24289 => "01101000", 24290 => "10101110", 24291 => "10100001", 24293 => "00101011", 24295 => "00011111", 24298 => "00100101", 24301 => "11101010", 24302 => "10100010", 24303 => "01001011", 24304 => "01000011", 24309 => "10111110", 24312 => "00000001", 24313 => "10101000", 24314 => "00011001", 24315 => "10100100", 24316 => "10111000", 24319 => "01000111", 24320 => "00001110", 24321 => "11001100", 24324 => "11011011", 24327 => "00111111", 24328 => "11111101", 24330 => "01110100", 24331 => "10101110", 24332 => "10011011", 24334 => "10110001", 24335 => "00001110", 24336 => "10010110", 24337 => "00001110", 24338 => "01100000", 24346 => "10011101", 24347 => "01011111", 24348 => "10111101", 24353 => "11000010", 24354 => "10101110", 24355 => "00001110", 24357 => "01001000", 24359 => "11000010", 24363 => "00111000", 24364 => "01001101", 24365 => "01011101", 24366 => "00110110", 24367 => "11100101", 24369 => "10010010", 24372 => "11110011", 24375 => "00010010", 24376 => "10011001", 24377 => "00000101", 24378 => "11100100", 24379 => "10000111", 24381 => "11111001", 24382 => "01110000", 24383 => "11101010", 24388 => "10100100", 24390 => "11011100", 24391 => "01001011", 24396 => "11000011", 24400 => "00111111", 24402 => "10010100", 24405 => "00011100", 24408 => "01010000", 24412 => "11100110", 24413 => "11100110", 24418 => "00001011", 24420 => "11111111", 24423 => "11011010", 24424 => "10100110", 24425 => "11110011", 24427 => "00101011", 24433 => "11101011", 24434 => "10001010", 24437 => "10110110", 24438 => "01001100", 24439 => "01001000", 24440 => "01100001", 24443 => "00010101", 24447 => "00010110", 24449 => "11100001", 24450 => "00101110", 24451 => "10101101", 24452 => "10010110", 24453 => "00101011", 24455 => "11110111", 24458 => "10011111", 24459 => "00011111", 24462 => "01101011", 24463 => "00111110", 24464 => "11011101", 24466 => "00000011", 24468 => "01000011", 24469 => "00011101", 24471 => "00100101", 24472 => "11111001", 24475 => "00111111", 24476 => "00010001", 24478 => "11000000", 24479 => "01011010", 24482 => "00110011", 24483 => "11010011", 24484 => "10100101", 24485 => "00101110", 24487 => "01010101", 24489 => "00111010", 24491 => "00000110", 24494 => "11000011", 24498 => "01011000", 24501 => "01001111", 24507 => "01111010", 24513 => "10111000", 24515 => "11000000", 24516 => "00011010", 24518 => "11110011", 24519 => "11010000", 24520 => "11000111", 24524 => "00100001", 24525 => "01001110", 24526 => "10010100", 24527 => "11110101", 24530 => "01011111", 24531 => "11101100", 24532 => "01001111", 24533 => "10001100", 24534 => "01011001", 24536 => "00101000", 24540 => "00001001", 24543 => "01110011", 24556 => "01111111", 24557 => "01101001", 24561 => "11001011", 24562 => "00110111", 24563 => "10000101", 24564 => "10110100", 24565 => "01010110", 24566 => "11011000", 24568 => "11000111", 24569 => "00010111", 24573 => "01001000", 24574 => "01001000", 24575 => "11111010", 24576 => "00000101", 24580 => "00010010", 24583 => "11101000", 24584 => "11110110", 24585 => "11011001", 24586 => "00010010", 24587 => "01110001", 24590 => "10000010", 24592 => "11111011", 24595 => "11110100", 24598 => "01100100", 24599 => "00111000", 24601 => "01001011", 24602 => "01010001", 24603 => "10101000", 24604 => "10011111", 24606 => "00011001", 24608 => "10001001", 24611 => "01000000", 24612 => "11010111", 24613 => "11010000", 24614 => "11101011", 24615 => "10110011", 24616 => "01001001", 24617 => "01000111", 24622 => "00000010", 24624 => "10000110", 24627 => "00010100", 24629 => "11001100", 24630 => "10010000", 24634 => "11110001", 24635 => "01100110", 24636 => "11001011", 24637 => "01111101", 24641 => "00001110", 24642 => "11001001", 24643 => "00011101", 24645 => "01101010", 24647 => "10011111", 24648 => "01101111", 24649 => "00111001", 24651 => "10100110", 24652 => "10001000", 24653 => "10100000", 24657 => "10110100", 24660 => "01111100", 24663 => "11111101", 24664 => "11110111", 24665 => "11000111", 24666 => "00010010", 24668 => "01110100", 24669 => "10110001", 24670 => "10010101", 24671 => "10010011", 24673 => "10000101", 24675 => "10001011", 24676 => "11110110", 24679 => "10001011", 24681 => "11111100", 24682 => "01101011", 24683 => "10000111", 24684 => "11011100", 24687 => "11010111", 24688 => "11110011", 24689 => "10000010", 24690 => "11001100", 24694 => "00011000", 24697 => "01111100", 24698 => "10000100", 24699 => "00001100", 24700 => "01111000", 24701 => "00011111", 24702 => "10101011", 24706 => "11110111", 24709 => "10000111", 24721 => "01111011", 24722 => "10101001", 24724 => "01110101", 24725 => "11110111", 24726 => "10001000", 24729 => "10111001", 24730 => "10010101", 24732 => "10101110", 24738 => "01010001", 24740 => "00011101", 24742 => "01011101", 24743 => "00010110", 24744 => "01111101", 24746 => "01110000", 24749 => "11010101", 24750 => "11110000", 24753 => "01011111", 24754 => "11000101", 24756 => "11010001", 24759 => "01000011", 24765 => "10101100", 24767 => "10100001", 24768 => "01111101", 24771 => "01101011", 24772 => "01001000", 24774 => "00101011", 24776 => "00100100", 24778 => "00111010", 24779 => "01110001", 24781 => "10000010", 24783 => "10111101", 24785 => "01011100", 24787 => "11110011", 24790 => "11011000", 24791 => "01110100", 24792 => "01110100", 24795 => "11101010", 24797 => "11000001", 24798 => "00111100", 24799 => "11000110", 24801 => "10111010", 24803 => "01000101", 24806 => "01010000", 24807 => "00100010", 24815 => "01110001", 24817 => "00110010", 24819 => "01001011", 24820 => "10110101", 24821 => "11011110", 24822 => "10001001", 24823 => "00100011", 24827 => "10110111", 24828 => "11000000", 24829 => "00011110", 24830 => "00001011", 24831 => "00001110", 24836 => "01101001", 24837 => "00001111", 24838 => "10100100", 24841 => "01011011", 24843 => "00001001", 24845 => "01011010", 24849 => "00010011", 24857 => "01110010", 24859 => "11111001", 24860 => "10110001", 24863 => "11011001", 24868 => "01111111", 24869 => "00001001", 24870 => "00101001", 24872 => "11001000", 24873 => "10111001", 24876 => "01101010", 24878 => "11101000", 24880 => "00111111", 24881 => "01110000", 24882 => "01001011", 24883 => "00011001", 24886 => "11001110", 24887 => "00110011", 24891 => "01110011", 24892 => "01011110", 24895 => "01100110", 24896 => "11011101", 24897 => "10111001", 24898 => "10100110", 24902 => "00101100", 24903 => "00001000", 24905 => "10111011", 24907 => "10111111", 24910 => "10011010", 24911 => "00001011", 24912 => "00101011", 24913 => "10011101", 24917 => "11110110", 24918 => "00010100", 24919 => "01010001", 24921 => "00011001", 24924 => "01010010", 24926 => "00110101", 24929 => "01000010", 24931 => "10011001", 24934 => "11100010", 24935 => "00000110", 24936 => "00110110", 24938 => "00111111", 24939 => "11110010", 24941 => "00011110", 24943 => "00111001", 24945 => "10001001", 24946 => "10101010", 24947 => "01101111", 24948 => "11011000", 24949 => "10110000", 24951 => "11110000", 24960 => "00111011", 24962 => "01111010", 24963 => "10100111", 24964 => "00001010", 24968 => "00011000", 24969 => "00100100", 24970 => "11001100", 24971 => "11010110", 24975 => "00011110", 24977 => "11011001", 24983 => "01000011", 24984 => "10110100", 24988 => "10101100", 24989 => "10110010", 24995 => "10111110", 25000 => "11000001", 25001 => "10110110", 25002 => "01000100", 25006 => "10111111", 25007 => "10101100", 25008 => "10111110", 25009 => "01110001", 25010 => "01101111", 25011 => "00101010", 25013 => "11011100", 25014 => "01100100", 25017 => "10001001", 25018 => "11011001", 25020 => "00101101", 25022 => "00110111", 25026 => "00110011", 25029 => "00000001", 25030 => "01001000", 25031 => "10110001", 25032 => "01110011", 25033 => "11011001", 25034 => "10111100", 25038 => "10000110", 25039 => "00000011", 25042 => "11100010", 25044 => "11111111", 25045 => "10111011", 25046 => "00001010", 25048 => "01010100", 25049 => "00000011", 25052 => "00101101", 25053 => "11001101", 25056 => "01000110", 25057 => "10101110", 25061 => "00111010", 25062 => "10000110", 25064 => "11011000", 25065 => "01001110", 25068 => "01001101", 25069 => "00010011", 25072 => "11001010", 25078 => "11011000", 25081 => "11101011", 25082 => "01100110", 25083 => "01110000", 25088 => "11100011", 25090 => "10000111", 25093 => "11110001", 25094 => "10001010", 25096 => "11000011", 25097 => "10010001", 25098 => "01100010", 25099 => "10011001", 25100 => "11101011", 25102 => "00000111", 25108 => "00010101", 25109 => "11010100", 25111 => "10100110", 25112 => "00101010", 25116 => "01001100", 25117 => "01011111", 25119 => "11000110", 25122 => "00000100", 25123 => "10110100", 25124 => "01011011", 25127 => "00010001", 25131 => "01001001", 25133 => "10111110", 25135 => "11110010", 25136 => "11101011", 25138 => "01100101", 25139 => "01000110", 25140 => "00100000", 25143 => "01001110", 25144 => "10010001", 25145 => "01001110", 25146 => "10011001", 25147 => "11110111", 25148 => "01001001", 25149 => "11100001", 25150 => "11001111", 25151 => "11100100", 25153 => "11011010", 25155 => "01010011", 25156 => "10011101", 25157 => "00100010", 25160 => "11100011", 25164 => "00111011", 25167 => "01110111", 25170 => "01011000", 25171 => "11001111", 25172 => "01101100", 25175 => "01111111", 25176 => "01110000", 25179 => "11111000", 25180 => "11001100", 25181 => "00011010", 25185 => "01100010", 25188 => "01010111", 25190 => "00001001", 25191 => "11110111", 25193 => "10100110", 25195 => "00011111", 25196 => "01000110", 25200 => "01110101", 25202 => "01110110", 25203 => "00111010", 25204 => "10100101", 25205 => "00000111", 25206 => "00010010", 25207 => "00011011", 25208 => "10111110", 25210 => "10101011", 25211 => "00110100", 25212 => "11101111", 25213 => "10011110", 25215 => "10000110", 25222 => "01001010", 25224 => "01101111", 25225 => "00010001", 25227 => "11110110", 25230 => "10111001", 25232 => "10010001", 25235 => "10111010", 25236 => "10100010", 25237 => "11110010", 25240 => "11111010", 25241 => "00100111", 25243 => "01101111", 25248 => "10000001", 25251 => "01000001", 25253 => "10001001", 25254 => "00111000", 25264 => "11001001", 25265 => "01011100", 25266 => "01110101", 25267 => "01100110", 25268 => "01111010", 25271 => "01001100", 25272 => "00101111", 25274 => "11010001", 25279 => "00001011", 25282 => "01011001", 25284 => "11111111", 25285 => "00100111", 25287 => "10101010", 25288 => "10001100", 25289 => "10010111", 25291 => "10110101", 25292 => "10010011", 25300 => "00100000", 25302 => "01010000", 25305 => "00111111", 25306 => "01010010", 25307 => "01001111", 25312 => "10001100", 25314 => "01111010", 25315 => "10010000", 25316 => "10111001", 25318 => "10001111", 25319 => "01111001", 25322 => "00010001", 25325 => "01010110", 25327 => "11101010", 25328 => "01111000", 25332 => "01000110", 25333 => "11001111", 25334 => "10111001", 25337 => "00001111", 25338 => "00000101", 25339 => "10000100", 25340 => "11001000", 25344 => "01111001", 25346 => "10110110", 25347 => "10000011", 25349 => "11011100", 25351 => "11010110", 25354 => "01011111", 25355 => "01001011", 25356 => "10111110", 25357 => "11010001", 25358 => "10010000", 25359 => "00010111", 25361 => "10010011", 25366 => "11010011", 25367 => "01000000", 25368 => "01001100", 25369 => "11010111", 25373 => "11101011", 25374 => "00010101", 25375 => "11101111", 25377 => "11110000", 25382 => "11100101", 25383 => "11100001", 25385 => "10011101", 25387 => "01110010", 25388 => "01100101", 25389 => "11000110", 25390 => "01101011", 25392 => "10100111", 25396 => "00000101", 25397 => "11010000", 25401 => "11100000", 25404 => "00110000", 25405 => "11010000", 25406 => "01000100", 25407 => "10111001", 25408 => "10100110", 25411 => "00101010", 25414 => "10100101", 25415 => "10110111", 25418 => "11001010", 25420 => "00000001", 25421 => "10111110", 25422 => "10000110", 25424 => "00001111", 25425 => "01110011", 25426 => "01111110", 25427 => "01000100", 25428 => "01110001", 25431 => "00011110", 25432 => "11111111", 25433 => "11110001", 25435 => "00110100", 25436 => "00011001", 25437 => "10110010", 25438 => "11101010", 25440 => "01010101", 25445 => "10110100", 25448 => "00001000", 25451 => "01000011", 25453 => "10100001", 25454 => "01010001", 25457 => "11100100", 25458 => "00110001", 25459 => "10101000", 25462 => "11111110", 25463 => "01101110", 25464 => "11111011", 25467 => "10110011", 25471 => "11100110", 25480 => "10100101", 25481 => "00110110", 25485 => "11001000", 25487 => "00010011", 25489 => "11111010", 25496 => "10110000", 25497 => "10101110", 25498 => "00001010", 25499 => "01001110", 25500 => "10001011", 25502 => "11101011", 25503 => "01100001", 25504 => "01001101", 25506 => "01010000", 25507 => "11101100", 25508 => "10100101", 25512 => "11011101", 25514 => "01010001", 25516 => "11101111", 25517 => "00101000", 25520 => "00101000", 25521 => "00001001", 25525 => "11110110", 25527 => "10101011", 25528 => "10101011", 25533 => "11111101", 25538 => "00100100", 25539 => "10010100", 25540 => "11000111", 25541 => "11110011", 25547 => "11101110", 25548 => "01101100", 25549 => "11010011", 25550 => "10100001", 25554 => "11011101", 25557 => "00100001", 25558 => "01101001", 25564 => "10100100", 25568 => "10010001", 25570 => "00011101", 25572 => "10101100", 25575 => "10011111", 25576 => "10000111", 25579 => "00001110", 25581 => "11111000", 25582 => "01110101", 25583 => "00000101", 25584 => "11000110", 25590 => "11000110", 25591 => "00000010", 25594 => "11001110", 25598 => "00011001", 25599 => "10111100", 25602 => "10100001", 25607 => "10000001", 25609 => "10110010", 25611 => "10101110", 25612 => "00000001", 25615 => "01000101", 25616 => "10011100", 25617 => "11001100", 25619 => "11101101", 25620 => "00011010", 25621 => "11000100", 25622 => "10001110", 25624 => "01001011", 25629 => "01111001", 25630 => "10101001", 25631 => "10001110", 25632 => "10100000", 25633 => "01011010", 25638 => "00010000", 25639 => "01001101", 25640 => "11000011", 25642 => "11000010", 25645 => "10001000", 25646 => "11010011", 25647 => "10011111", 25648 => "01111100", 25649 => "00111110", 25650 => "00010111", 25654 => "11011110", 25658 => "01111000", 25659 => "11101111", 25660 => "01100101", 25661 => "01110101", 25662 => "00010100", 25666 => "00101000", 25668 => "11001100", 25669 => "11101010", 25670 => "10111101", 25674 => "10010101", 25676 => "11111100", 25677 => "11000101", 25678 => "01111001", 25680 => "01010000", 25681 => "11010100", 25682 => "11010010", 25683 => "00011101", 25684 => "00000010", 25685 => "11110000", 25687 => "10001001", 25688 => "00100110", 25689 => "00001101", 25692 => "10011000", 25693 => "01100000", 25694 => "11111101", 25699 => "01101111", 25700 => "10110100", 25704 => "11101110", 25705 => "00101000", 25708 => "11011101", 25709 => "11000000", 25710 => "00100010", 25716 => "01011010", 25719 => "00101010", 25720 => "10111000", 25724 => "10100001", 25726 => "10100000", 25727 => "01011010", 25728 => "00100100", 25729 => "10010001", 25731 => "10011110", 25737 => "01111111", 25742 => "11111010", 25743 => "01110111", 25750 => "11111101", 25754 => "00011011", 25756 => "11110100", 25760 => "00111000", 25763 => "01111101", 25767 => "11100000", 25768 => "01111110", 25769 => "01110100", 25771 => "00110001", 25776 => "00001000", 25778 => "10011110", 25780 => "01101011", 25781 => "11110000", 25784 => "01111101", 25788 => "00101010", 25791 => "10000001", 25792 => "11011101", 25793 => "10001110", 25794 => "01001000", 25795 => "10101000", 25797 => "11001101", 25798 => "00100100", 25799 => "01001011", 25802 => "11101011", 25803 => "10001010", 25804 => "01011111", 25808 => "11001101", 25809 => "10010001", 25810 => "10000101", 25816 => "01111100", 25818 => "10000100", 25819 => "00101000", 25822 => "01001011", 25824 => "11101000", 25828 => "01001111", 25831 => "00011100", 25832 => "01001110", 25833 => "11011011", 25835 => "11110110", 25836 => "11111110", 25837 => "01010001", 25838 => "00100001", 25840 => "00100000", 25842 => "10111101", 25843 => "00110010", 25845 => "00001011", 25846 => "00011011", 25849 => "11011000", 25850 => "11011100", 25851 => "10110110", 25852 => "11101001", 25854 => "01010110", 25860 => "00111010", 25861 => "01110111", 25863 => "01001010", 25865 => "01011010", 25866 => "00110110", 25867 => "10011100", 25869 => "10000100", 25870 => "10100111", 25873 => "11001010", 25875 => "00110011", 25876 => "10010010", 25877 => "01100101", 25878 => "01001000", 25879 => "01011010", 25883 => "10000110", 25885 => "01101000", 25888 => "01101010", 25889 => "11111000", 25891 => "01010100", 25894 => "11100111", 25895 => "01011001", 25896 => "00110001", 25899 => "01000011", 25900 => "10111010", 25901 => "11000110", 25902 => "01011101", 25904 => "11000111", 25905 => "11110110", 25906 => "01000001", 25907 => "10000000", 25908 => "00011111", 25909 => "10011110", 25911 => "00101101", 25912 => "11000010", 25913 => "10010101", 25920 => "01100110", 25921 => "11011111", 25926 => "11011010", 25927 => "01100110", 25928 => "10100001", 25929 => "00110111", 25931 => "10101001", 25933 => "10001001", 25936 => "10110101", 25938 => "11010011", 25940 => "11101011", 25941 => "10101010", 25943 => "11100001", 25944 => "00001110", 25947 => "10111111", 25952 => "10001110", 25955 => "01011000", 25958 => "11101001", 25959 => "00000100", 25963 => "10110100", 25964 => "10000010", 25965 => "11000011", 25966 => "00100101", 25967 => "00011100", 25968 => "01100110", 25970 => "01011100", 25972 => "00011101", 25974 => "00101110", 25975 => "10001010", 25979 => "10000001", 25980 => "10001101", 25981 => "11100010", 25984 => "10111111", 25985 => "00100001", 25986 => "01101000", 25987 => "11001111", 25988 => "11100110", 25990 => "01010011", 25991 => "11000111", 25994 => "10011001", 25995 => "10100000", 25996 => "11110110", 25998 => "01101010", 26000 => "11101101", 26002 => "00010100", 26003 => "00100101", 26005 => "01001111", 26006 => "01101000", 26007 => "11000011", 26009 => "00111000", 26010 => "11000111", 26011 => "01000010", 26012 => "10010101", 26013 => "01101111", 26014 => "01110010", 26016 => "10000001", 26018 => "00100110", 26019 => "11001010", 26020 => "11110010", 26021 => "00010010", 26022 => "11100011", 26023 => "00111000", 26027 => "10111000", 26030 => "11010101", 26033 => "01011101", 26034 => "00100001", 26036 => "00000101", 26037 => "10110110", 26038 => "11100111", 26041 => "01100101", 26042 => "10001110", 26044 => "11000100", 26045 => "00111001", 26049 => "10010011", 26051 => "11010001", 26052 => "00101010", 26058 => "11001010", 26062 => "11100110", 26066 => "01101001", 26067 => "11001101", 26070 => "11110111", 26072 => "10011110", 26073 => "10010110", 26074 => "00101011", 26076 => "01001110", 26078 => "00101010", 26080 => "00010001", 26081 => "00111001", 26084 => "10001111", 26086 => "11001001", 26087 => "10010100", 26088 => "01101111", 26089 => "11101101", 26093 => "00111011", 26094 => "11001100", 26095 => "11111110", 26100 => "10010100", 26102 => "11000111", 26104 => "11011111", 26105 => "01111100", 26107 => "11011000", 26109 => "01011111", 26110 => "10110001", 26111 => "10000111", 26112 => "11000000", 26113 => "10101001", 26114 => "01000011", 26118 => "11010000", 26124 => "01101001", 26125 => "00100001", 26127 => "10110100", 26128 => "01111011", 26130 => "01100110", 26132 => "00110110", 26136 => "00011111", 26139 => "10011111", 26143 => "01000001", 26145 => "01001101", 26150 => "11100000", 26151 => "11101110", 26157 => "00111001", 26158 => "11011111", 26159 => "01100010", 26160 => "11010000", 26162 => "10010100", 26163 => "00110111", 26164 => "10000001", 26167 => "11011000", 26168 => "11010111", 26171 => "11100111", 26172 => "11111000", 26173 => "10011011", 26174 => "10110111", 26176 => "00010101", 26177 => "10110101", 26181 => "01101100", 26182 => "01110000", 26183 => "01100001", 26184 => "01000111", 26187 => "01101100", 26188 => "00011101", 26189 => "00000001", 26196 => "01011100", 26197 => "11100110", 26199 => "01100100", 26200 => "01011110", 26201 => "11111011", 26202 => "01010010", 26204 => "10101000", 26207 => "00011010", 26208 => "11101111", 26210 => "10100100", 26211 => "01110011", 26214 => "00000100", 26217 => "11100010", 26219 => "00001010", 26220 => "10011111", 26221 => "11110000", 26222 => "01000101", 26224 => "01001001", 26227 => "00101100", 26228 => "11111000", 26230 => "00001100", 26231 => "11100001", 26232 => "10000111", 26235 => "00011010", 26237 => "01010001", 26242 => "01100110", 26243 => "00010001", 26246 => "11011110", 26249 => "00000011", 26251 => "00001111", 26252 => "10100011", 26259 => "11101001", 26261 => "00010100", 26264 => "00010011", 26265 => "00011010", 26269 => "01111110", 26270 => "11111010", 26272 => "00011000", 26274 => "00010111", 26288 => "10100010", 26289 => "01001110", 26290 => "11000011", 26292 => "10010100", 26293 => "01011010", 26294 => "11011100", 26295 => "11011011", 26297 => "11111110", 26298 => "01001001", 26303 => "00100110", 26306 => "00001100", 26308 => "10110100", 26310 => "10111011", 26312 => "01101111", 26317 => "11100111", 26318 => "01000000", 26319 => "01001101", 26321 => "00010000", 26325 => "11011010", 26328 => "10011000", 26329 => "01010011", 26334 => "01000011", 26341 => "10110011", 26342 => "11000110", 26343 => "00010100", 26344 => "11010001", 26345 => "11001011", 26346 => "10001010", 26348 => "10111001", 26350 => "01000100", 26351 => "00000100", 26352 => "00001111", 26354 => "10101011", 26355 => "01111011", 26357 => "10100001", 26360 => "01010011", 26361 => "11000101", 26362 => "10100001", 26367 => "10011001", 26368 => "00001110", 26369 => "10011110", 26370 => "11100011", 26374 => "01110101", 26376 => "00100011", 26379 => "01111101", 26383 => "11100111", 26384 => "01001010", 26387 => "11100110", 26388 => "11110100", 26391 => "00011001", 26392 => "00001001", 26393 => "01000000", 26395 => "11011001", 26398 => "11010110", 26399 => "01101000", 26401 => "11010100", 26403 => "00001000", 26407 => "01111111", 26409 => "10001010", 26413 => "11000010", 26414 => "00101101", 26415 => "11100001", 26417 => "10001100", 26420 => "01111110", 26421 => "00101001", 26424 => "10111101", 26425 => "10011010", 26426 => "10100111", 26429 => "11100111", 26432 => "01011101", 26433 => "00000111", 26434 => "00001001", 26435 => "11000001", 26436 => "11001011", 26438 => "10001100", 26439 => "01011100", 26440 => "11010111", 26441 => "11011010", 26445 => "11011001", 26451 => "01000001", 26453 => "10100111", 26454 => "10010100", 26457 => "11011111", 26461 => "01000001", 26470 => "01011101", 26471 => "00001011", 26477 => "10001110", 26478 => "10111011", 26479 => "00011111", 26480 => "11001111", 26481 => "01111000", 26482 => "00001100", 26485 => "11101100", 26486 => "01100011", 26487 => "10011000", 26488 => "00010011", 26490 => "01100111", 26491 => "11100111", 26493 => "01110001", 26494 => "01101000", 26495 => "00101111", 26496 => "11011000", 26498 => "10111111", 26502 => "01000011", 26503 => "11011100", 26505 => "00001100", 26507 => "01011110", 26508 => "00001001", 26509 => "10010110", 26510 => "00100001", 26511 => "01100011", 26514 => "10110111", 26515 => "00001011", 26517 => "00011110", 26518 => "00101110", 26524 => "11111110", 26526 => "01101010", 26529 => "01011010", 26530 => "00101101", 26531 => "10001110", 26532 => "01000110", 26535 => "00000011", 26537 => "01011101", 26539 => "11011100", 26541 => "10111010", 26542 => "10101110", 26547 => "10000101", 26551 => "10100011", 26555 => "11010011", 26557 => "10010000", 26558 => "11111100", 26560 => "11001110", 26561 => "01111010", 26562 => "00100110", 26564 => "10111111", 26565 => "01000001", 26566 => "10101100", 26568 => "10111110", 26570 => "11011010", 26577 => "10101001", 26579 => "10110110", 26580 => "01100011", 26583 => "10101010", 26585 => "10101100", 26586 => "01000100", 26589 => "01110011", 26590 => "00100001", 26591 => "01011001", 26592 => "11010110", 26594 => "01011010", 26595 => "01001001", 26596 => "01001011", 26597 => "01111101", 26598 => "11011111", 26600 => "10111010", 26606 => "11010110", 26608 => "10110011", 26611 => "10101111", 26612 => "00011110", 26614 => "01010011", 26615 => "01110101", 26619 => "00110101", 26620 => "11100010", 26621 => "11111111", 26622 => "10010011", 26623 => "10110000", 26626 => "11001011", 26627 => "01010000", 26628 => "10110100", 26631 => "00001011", 26632 => "01111100", 26633 => "01100011", 26635 => "10111011", 26637 => "01101010", 26639 => "01000010", 26640 => "10001110", 26641 => "01010001", 26642 => "10010110", 26643 => "11101101", 26644 => "01011001", 26647 => "01111010", 26649 => "10100100", 26650 => "01101011", 26652 => "01010010", 26654 => "01111001", 26659 => "01010010", 26660 => "11011011", 26661 => "01110000", 26663 => "11111111", 26664 => "10111000", 26666 => "00111011", 26667 => "10011011", 26670 => "00100110", 26672 => "11011001", 26673 => "10110001", 26675 => "11101101", 26677 => "01111100", 26678 => "01111100", 26681 => "01110001", 26682 => "01010101", 26684 => "10010000", 26685 => "01111101", 26686 => "10010011", 26687 => "01010110", 26690 => "11000101", 26691 => "00000101", 26692 => "00000001", 26693 => "00111000", 26696 => "00111010", 26697 => "10111100", 26698 => "00101101", 26703 => "10000110", 26704 => "11100110", 26706 => "10010010", 26707 => "10010100", 26709 => "10011000", 26710 => "11100111", 26712 => "10111001", 26716 => "11100001", 26717 => "10001001", 26720 => "01110100", 26721 => "10011001", 26722 => "11101111", 26723 => "01011110", 26724 => "10011111", 26725 => "00001111", 26727 => "11010100", 26729 => "10001011", 26730 => "01100101", 26731 => "01111110", 26733 => "00111001", 26735 => "11000111", 26738 => "01000110", 26739 => "00111110", 26740 => "10010100", 26741 => "10101101", 26746 => "10000111", 26748 => "00010110", 26749 => "01011000", 26752 => "11101010", 26753 => "01100010", 26755 => "01110110", 26756 => "01100001", 26758 => "11010100", 26759 => "11010001", 26762 => "00011111", 26763 => "00011000", 26765 => "00011110", 26767 => "00010100", 26768 => "11010110", 26769 => "01111110", 26774 => "10100100", 26775 => "01101101", 26777 => "00101010", 26779 => "11101111", 26785 => "10101010", 26786 => "11111101", 26787 => "01011111", 26792 => "00110000", 26794 => "11111011", 26795 => "11011011", 26796 => "11111110", 26797 => "10100100", 26799 => "00111100", 26800 => "11111001", 26802 => "00110111", 26803 => "00100010", 26805 => "00010100", 26808 => "10000100", 26811 => "00110110", 26813 => "10001100", 26817 => "00000111", 26818 => "11001100", 26820 => "10111000", 26821 => "00100100", 26822 => "11011101", 26823 => "10000111", 26824 => "01011001", 26827 => "01110111", 26829 => "01001100", 26833 => "01101011", 26834 => "01011101", 26835 => "01110110", 26836 => "01000100", 26838 => "10110101", 26839 => "01001011", 26844 => "01100111", 26851 => "00001010", 26853 => "10110111", 26854 => "01101101", 26855 => "10110010", 26857 => "11101000", 26859 => "01100110", 26861 => "10011101", 26863 => "11000001", 26864 => "01111111", 26867 => "01000111", 26868 => "01000111", 26869 => "01010000", 26870 => "11111011", 26873 => "01001000", 26874 => "00111100", 26875 => "01101011", 26877 => "10011001", 26878 => "11101001", 26880 => "11001111", 26881 => "11010100", 26882 => "10100001", 26883 => "01110110", 26884 => "01101111", 26887 => "00000011", 26890 => "11110001", 26892 => "10100001", 26893 => "11010001", 26895 => "10110100", 26898 => "00100100", 26901 => "11000001", 26903 => "10111111", 26904 => "11011000", 26905 => "11000111", 26909 => "00001011", others => (others =>'0'));component project_reti_logiche is 
    port (
            i_clk         : in  std_logic;
            i_start       : in  std_logic;
            i_rst         : in  std_logic;
            i_data       : in  std_logic_vector(7 downto 0); --1 byte
            o_address     : out std_logic_vector(15 downto 0); --16 bit addr: max size is 255*255 + 3 more for max x and y and thresh.
            o_done            : out std_logic;
            o_en         : out std_logic;
            o_we       : out std_logic;
            o_data            : out std_logic_vector (7 downto 0)
          );
end component project_reti_logiche;


begin 
	UUT: project_reti_logiche
	port map (
		  i_clk      	=> tb_clk,	
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address, 
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
		  o_we 	=> mem_we,
          o_data    => mem_i_data
);

p_CLK_GEN : process is
  begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
  end process p_CLK_GEN; 
  
  
MEM : process(tb_clk)
   begin
    if tb_clk'event and tb_clk = '1' then
     if enable_wire = '1' then
      if mem_we = '1' then
       RAM(conv_integer(mem_address))              <= mem_i_data;
       mem_o_data                      <= mem_i_data after 1 ns;
      else
       mem_o_data <= RAM(conv_integer(mem_address)) after 1 ns;
      end if;
     end if;
    end if;
   end process;
 
  
test : process is
begin 
wait for 100 ns;
wait for c_CLOCK_PERIOD;
tb_rst <= '1';
wait for c_CLOCK_PERIOD;
tb_rst <= '0';
wait for c_CLOCK_PERIOD;
tb_start <= '1';
wait for c_CLOCK_PERIOD; 
tb_start <= '0';
wait until tb_done = '1';
wait until tb_done = '0';
wait until rising_edge(tb_clk); 

assert RAM(1) = "01101001" report "FAIL high bits" severity failure;
assert RAM(0) = "00011110" report "FAIL low bits" severity failure;
assert false report "Simulation Ended!, test passed" severity failure;
end process test;
end projecttb;