----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 12.12.2017 17:48:44
-- Design Name: 
-- Module Name: FSM_testbench - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
 
entity project_tb is
end project_tb;


architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 15 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst		    : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		    : std_logic := '0';
signal   mem_o_data,mem_i_data		: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		: std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (2 => "01001110", 3 => "00010010", 4 => "01000100", 8 => "11101111", 12 => "11001011", 13 => "01000001", 16 => "01110000", 18 => "10100010", 19 => "00011001", 20 => "01001001", 25 => "11110111", 26 => "00011111", 28 => "01011010", 33 => "10110110", 34 => "00010111", 35 => "00000110", 36 => "10010110", 43 => "11000100", 45 => "01111000", 46 => "00111101", 59 => "00111001", 65 => "11100111", 69 => "10000110", 70 => "00100000", 73 => "10010110", 74 => "11000100", 77 => "10010110", 78 => "11100111", 80 => "10001111", 85 => "01110011", 86 => "01111101", 91 => "11001000", 92 => "01101101", 94 => "00111011", 96 => "11110100", 97 => "11000001", 103 => "00001011", 106 => "11001000", 109 => "00101010", 110 => "10100010", 113 => "01001101", 115 => "01110010", 116 => "01100000", 122 => "11001000", 126 => "10011101", 135 => "01111000", 145 => "11101010", 149 => "10110110", 150 => "11011110", 153 => "11101110", 156 => "00110100", 158 => "10101010", 160 => "11001110", 162 => "00011101", 172 => "01011010", 178 => "00000111", 180 => "01110111", 181 => "10111000", 182 => "11110101", 183 => "10001010", 186 => "11110001", 191 => "10001000", 193 => "01100001", 196 => "01101011", 197 => "00111011", 200 => "10010010", 204 => "10110011", 206 => "11110010", 207 => "10011111", 210 => "10111010", 215 => "00110010", 224 => "01000110", 233 => "01001110", 239 => "00111001", 241 => "10101001", 244 => "10010100", 245 => "00110101", 247 => "00111101", 251 => "00001000", 252 => "10111110", 253 => "10111110", 262 => "00011101", 266 => "00110010", 267 => "01010011", 273 => "00010111", 274 => "00111101", 283 => "11110010", 284 => "10111011", 297 => "01001101", 301 => "00001111", 305 => "00101011", 306 => "00010011", 307 => "10111110", 310 => "10011100", 311 => "01010010", 316 => "10100101", 319 => "10100111", 320 => "01011010", 327 => "10101110", 328 => "00110111", 332 => "01001101", 333 => "11100110", 334 => "00011110", 335 => "11101001", 337 => "00001101", 339 => "10001000", 340 => "11000011", 341 => "01010011", 342 => "10000000", 345 => "11001110", 347 => "01111001", 350 => "11100011", 352 => "10001001", 356 => "11110110", 361 => "11100100", 363 => "01101010", 364 => "11000010", 375 => "11111001", 391 => "01010110", 392 => "01000100", 396 => "00110111", 398 => "11011011", 401 => "11011000", 402 => "10010111", 403 => "11010110", 405 => "01110010", 406 => "10100101", 413 => "01010010", 415 => "01110110", 416 => "11101100", 417 => "01011000", 419 => "10011101", 423 => "11001001", 425 => "11001000", 435 => "00001001", 437 => "01111110", 443 => "11000101", 444 => "00000010", 446 => "01110101", 452 => "11001100", 456 => "01111011", 457 => "01101111", 464 => "00011011", 466 => "10010000", 468 => "11100001", 470 => "00110111", 472 => "11000000", 475 => "00000111", 477 => "11011100", 485 => "11011010", 489 => "00101101", 490 => "00100111", 493 => "10011011", 494 => "11001000", 496 => "00111101", 498 => "01000101", 499 => "01100010", 503 => "10000011", 505 => "11110100", 507 => "01100000", 509 => "01000000", 512 => "01100110", 514 => "00010111", 520 => "00101100", 529 => "01100000", 531 => "10100110", 533 => "00111101", 535 => "01100101", 536 => "11011100", 539 => "10110011", 542 => "10000001", 546 => "10100110", 548 => "00111110", 552 => "00101100", 555 => "01110100", 561 => "00110110", 564 => "00110001", 565 => "01000010", 566 => "01000010", 569 => "10111000", 573 => "10001010", 579 => "01000011", 586 => "10100110", 589 => "10110001", 593 => "01011011", 595 => "11010101", 596 => "01000001", 600 => "01100010", 603 => "01010010", 604 => "10101001", 607 => "01101101", 611 => "00100000", 612 => "01110111", 616 => "11101000", 617 => "10111010", 620 => "11011110", 621 => "01110100", 623 => "00100001", 624 => "11011101", 625 => "10010100", 628 => "11000101", 632 => "10001000", 638 => "10100101", 640 => "10011110", 642 => "01001100", 645 => "00001010", 647 => "00001011", 652 => "01100001", 665 => "11110010", 669 => "11011110", 671 => "11100010", 674 => "11101111", 676 => "10011110", 682 => "11000100", 683 => "10100100", 684 => "10010100", 687 => "10101100", 690 => "10100100", 691 => "01001000", 692 => "00001011", 693 => "01101110", 694 => "10000001", 700 => "00000111", 703 => "00110000", 706 => "01110001", 707 => "00100010", 708 => "00001001", 709 => "00100100", 710 => "00111011", 712 => "10100001", 717 => "01100001", 721 => "11110011", 726 => "11111110", 729 => "10100100", 731 => "10011011", 732 => "11110001", 733 => "01010000", 735 => "01001010", 736 => "10101110", 743 => "11111010", 744 => "11011001", 747 => "10001011", 755 => "01010000", 759 => "10101011", 765 => "00111111", 768 => "11111000", 772 => "10010010", 774 => "11111001", 775 => "00011001", 777 => "11100000", 778 => "11110100", 784 => "01100010", 789 => "10110010", 793 => "01111110", 795 => "00110010", 805 => "01111000", 807 => "10000110", 808 => "00101010", 809 => "01010000", 811 => "10011000", 813 => "01011000", 818 => "00110111", 822 => "11011101", 823 => "01110110", 829 => "11100001", 834 => "11011111", 835 => "00100110", 836 => "00010100", 837 => "00001011", 848 => "00111100", 851 => "00110000", 855 => "01010001", 861 => "11100101", 862 => "10010011", 867 => "11110100", 878 => "01101111", 882 => "01000011", 884 => "10110110", 886 => "10101111", 889 => "10101110", 894 => "11110100", 897 => "10111000", 899 => "01111001", 900 => "01011101", 902 => "00001110", 903 => "10101010", 905 => "11101000", 907 => "10001100", 909 => "00011010", 914 => "11111111", 923 => "00011000", 933 => "11010111", 935 => "00010100", 940 => "00010110", 941 => "11000111", 944 => "10000100", 946 => "01100100", 951 => "00101001", 952 => "00101110", 954 => "10000110", 962 => "11100001", 964 => "01110110", 966 => "11111111", 969 => "10001001", 970 => "10101111", 975 => "00000101", 981 => "10010000", 984 => "00110010", 985 => "00101110", 988 => "10101110", 990 => "01101010", 991 => "01110000", 992 => "11111111", 993 => "10011001", 994 => "10110101", 1001 => "10011111", 1002 => "00101110", 1003 => "01100001", 1009 => "00000111", 1011 => "00110000", 1015 => "00001100", 1017 => "10001110", 1020 => "01000101", 1022 => "01100110", 1024 => "01000010", 1031 => "01111000", 1034 => "10110011", 1036 => "00110010", 1045 => "11001100", 1047 => "00100001", 1051 => "00100100", 1054 => "10001101", 1062 => "10101100", 1065 => "10010110", 1066 => "00011010", 1068 => "01111000", 1071 => "00101110", 1073 => "10011010", 1075 => "00011100", 1077 => "01011011", 1078 => "01101011", 1081 => "01000011", 1083 => "01001001", 1093 => "00111010", 1099 => "10100111", 1100 => "10100000", 1105 => "00011110", 1124 => "11110111", 1126 => "11000110", 1128 => "00001010", 1130 => "11000010", 1132 => "10011101", 1138 => "00100111", 1140 => "01100010", 1141 => "00101000", 1158 => "10110110", 1159 => "10000111", 1160 => "00101011", 1161 => "01101001", 1163 => "01010000", 1164 => "00010111", 1165 => "00010001", 1167 => "11011101", 1168 => "01100101", 1169 => "01011101", 1172 => "01010101", 1174 => "11101001", 1178 => "00010100", 1179 => "11111000", 1180 => "10111011", 1187 => "01100000", 1193 => "10000101", 1194 => "01101001", 1203 => "00001010", 1206 => "01010010", 1207 => "01010110", 1211 => "01011011", 1212 => "10011101", 1216 => "11100110", 1218 => "01101111", 1220 => "00000110", 1224 => "01100010", 1230 => "01011111", 1231 => "01001010", 1234 => "00000001", 1238 => "11100011", 1241 => "00111010", 1243 => "01101101", 1245 => "01001110", 1247 => "10101011", 1258 => "11000001", 1261 => "01011001", 1262 => "11000111", 1267 => "11101001", 1271 => "01101111", 1273 => "01011101", 1278 => "01000111", 1281 => "11001111", 1282 => "10011101", 1284 => "10001101", 1286 => "10100101", 1289 => "10111110", 1291 => "00101100", 1294 => "01001001", 1295 => "10100001", 1301 => "10101100", 1305 => "00010101", 1319 => "10001101", 1326 => "10101111", 1329 => "11100010", 1334 => "11111111", 1335 => "11001010", 1336 => "01010110", 1341 => "01011011", 1344 => "01100001", 1345 => "00011011", 1348 => "10011000", 1349 => "00001100", 1355 => "01010011", 1356 => "01011010", 1357 => "00110000", 1361 => "11110001", 1368 => "00001011", 1369 => "10111001", 1373 => "10100001", 1374 => "00110011", 1375 => "00001100", 1378 => "11111111", 1381 => "00010100", 1387 => "10000001", 1390 => "00000101", 1391 => "00110001", 1392 => "01011110", 1393 => "11001101", 1396 => "00011100", 1398 => "01100110", 1400 => "11110001", 1401 => "00011100", 1403 => "01010100", others => (others =>'0'));component project_reti_logiche is 
    port (
            i_clk         : in  std_logic;
            i_start       : in  std_logic;
            i_rst         : in  std_logic;
            i_data       : in  std_logic_vector(7 downto 0); --1 byte
            o_address     : out std_logic_vector(15 downto 0); --16 bit addr: max size is 255*255 + 3 more for max x and y and thresh.
            o_done            : out std_logic;
            o_en         : out std_logic;
            o_we       : out std_logic;
            o_data            : out std_logic_vector (7 downto 0)
          );
end component project_reti_logiche;


begin 
	UUT: project_reti_logiche
	port map (
		  i_clk      	=> tb_clk,	
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address, 
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
		  o_we 	=> mem_we,
          o_data    => mem_i_data
);

p_CLK_GEN : process is
  begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
  end process p_CLK_GEN; 
  
  
MEM : process(tb_clk)
   begin
    if tb_clk'event and tb_clk = '1' then
     if enable_wire = '1' then
      if mem_we = '1' then
       RAM(conv_integer(mem_address))              <= mem_i_data;
       mem_o_data                      <= mem_i_data after 1 ns;
      else
       mem_o_data <= RAM(conv_integer(mem_address)) after 1 ns;
      end if;
     end if;
    end if;
   end process;
 
  
test : process is
begin 
wait for 100 ns;
wait for c_CLOCK_PERIOD;
tb_rst <= '1';
wait for c_CLOCK_PERIOD;
tb_rst <= '0';
wait for c_CLOCK_PERIOD;
tb_start <= '1';
wait for c_CLOCK_PERIOD; 
tb_start <= '0';
wait until tb_done = '1';
wait until tb_done = '0';
wait until rising_edge(tb_clk); 

assert RAM(1) = "00000101" report "FAIL high bits" severity failure;
assert RAM(0) = "01111100" report "FAIL low bits" severity failure;
assert false report "Simulation Ended!, test passed" severity failure;
end process test;
end projecttb;